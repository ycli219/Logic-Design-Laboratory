`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/12/04 14:32:25
// Design Name: 
// Module Name: lab7_2
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module clock_divider #(parameter n=25) (
    input clk,
    output reg clk_div
    );
    
    reg [31:0] count = 32'b0;
    always @(posedge clk) begin
        count <= count + 1'b1;
        if(count >= (2**n)-1) count <= 32'b0;
        clk_div <= (count < (2**n)/2) ? 1'b1 : 1'b0;
    end
endmodule


module lab7_2(
    input clk,
    input rst,
    input hold,
    inout PS2_CLK,
    inout PS2_DATA,
    output [3:0] vgaRed,
    output [3:0] vgaGreen,
    output [3:0] vgaBlue,
    output hsync,
    output vsync,
    output wire pass
    );
    
    wire de_hold;
    debounce m1(de_hold , hold , clk);
    
    
    parameter [8:0] LEFT_SHIFT_CODES  = 9'b0_0001_0010;
	parameter [8:0] RIGHT_SHIFT_CODES = 9'b0_0101_1001;
	parameter [8:0] KEY_CODES [0:11] = {
		9'b0_0100_0100,	// O => 44
		9'b0_0100_1101,	// P => 4D
		9'b0_0101_0100,	// [ => 54
		9'b0_0101_1011,	// ] => 5B
		9'b0_0100_0010,	// K => 42
		9'b0_0100_1011,	// L => 4B
		9'b0_0100_1100,	// ; => 4C
		9'b0_0101_0010,	// ' => 52
		9'b0_0011_1010,	// M => 3A
		9'b0_0100_0001,	// , => 41
		9'b0_0100_1001,  //. => 49
		9'b0_0100_1010   /// => 4A
	};
	
    wire [511:0] key_down;
	wire [8:0] last_change;
	wire been_ready;
	reg [3:0] key_num;
	
	
	KeyboardDecoder key_de (
		.key_down(key_down),
		.last_change(last_change),
		.key_valid(been_ready),
		.PS2_DATA(PS2_DATA),
		.PS2_CLK(PS2_CLK),
		.rst(rst),
		.clk(clk)
	);
	
	always @ (*) begin
		case (last_change)
			KEY_CODES[00] : key_num = 4'b0000;
			KEY_CODES[01] : key_num = 4'b0001;
			KEY_CODES[02] : key_num = 4'b0010;
			KEY_CODES[03] : key_num = 4'b0011;
			KEY_CODES[04] : key_num = 4'b0100;
			KEY_CODES[05] : key_num = 4'b0101;
			KEY_CODES[06] : key_num = 4'b0110;
			KEY_CODES[07] : key_num = 4'b0111;
			KEY_CODES[08] : key_num = 4'b1000;
			KEY_CODES[09] : key_num = 4'b1001;
			KEY_CODES[10] : key_num = 4'b1010;
			KEY_CODES[11] : key_num = 4'b1011;
			default: key_num = 4'b1111;
		endcase
	end
	
	
	wire shift;
	assign shift = (key_down[LEFT_SHIFT_CODES] == 1'b1 || key_down[RIGHT_SHIFT_CODES] == 1'b1) ? 1'b1 : 1'b0;
	
   reg [1:0] zero = 2'd0;
   reg [1:0] one = 2'd1;
   reg [1:0] two = 2'd2;
   reg [1:0] three = 2'd3;
   reg [1:0] four = 2'd3;
   reg [1:0] five = 2'd2;
   reg [1:0] six = 2'd1;
   reg [1:0] seven = 2'd0;
   reg [1:0] eight = 2'd1;
   reg [1:0] nine = 2'd0;
   reg [1:0] ten = 2'd3;
   reg [1:0] ele = 2'd2;
	
	
	//reg [3:0] rotate = 4'd13;
	always @(posedge clk or posedge rst) begin
	       if(rst == 1) begin
	           zero <= 2'd0;
               one <= 2'd1;
               two <= 2'd2;
               three <= 2'd3;
               four <= 2'd3;
               five <= 2'd2;
               six <= 2'd1;
               seven <= 2'd0;
               eight <= 2'd1;
               nine <= 2'd0;
               ten <= 2'd3;
               ele <= 2'd2;
	       end else begin
			if(been_ready && key_down[last_change] == 1'b1) begin
				if(key_num != 4'b1111 && pass == 0 && hold == 0) begin
					if(key_num == 4'd0) begin
                        if(shift == 1'b1) zero <= zero - 1;
                        else zero <= zero + 1;
                    end else if(key_num == 4'd1) begin
                        if(shift == 1'b1) one <= one - 1;
                        else one <= one + 1;
                    end else if(key_num == 4'd2) begin
                        if(shift == 1'b1) two <= two - 1;
                        else two <= two + 1;
                    end else if(key_num == 4'd3) begin
                        if(shift == 1'b1) three <= three - 1;
                        else three <= three + 1;
                    end else if(key_num == 4'd4) begin
                        if(shift == 1'b1) four <= four - 1;
                        else four <= four + 1;
                    end else if(key_num == 4'd5) begin
                        if(shift == 1'b1) five <= five - 1;
                        else five <= five + 1;
                    end else if(key_num == 4'd6) begin
                        if(shift == 1'b1) six <= six - 1;
                        else six <= six + 1;
                    end else if(key_num == 4'd7) begin
                        if(shift == 1'b1) seven <= seven - 1;
                        else seven <= seven + 1;
                    end else if(key_num == 4'd8) begin
                        if(shift == 1'b1) eight <= eight - 1;
                        else eight <= eight + 1;
                    end else if(key_num == 4'd9) begin
                        if(shift == 1'b1) nine <= nine - 1;
                        else nine <= nine + 1;
                    end else if(key_num == 4'd10) begin
                        if(shift == 1'b1) ten <= ten - 1;
                        else ten <= ten + 1;
                    end else if(key_num == 4'd11) begin
                        if(shift == 1'b1) ele <= ele - 1;
                        else ele <= ele + 1;
                    end
				end
			 end
			end
	end


    wire [11:0] data;
    wire clk_25MHz;
    reg [16:0] pixel_addr;
    wire [11:0] pixel;
    wire valid;
    wire [9:0] h_cnt;
    wire [9:0] v_cnt;
    
    clock_divider #(2) m2(clk,clk_25MHz);
    
    vga_controller vga_inst(
      .pclk(clk_25MHz),
      .reset(rst),
      .hsync(hsync),
      .vsync(vsync),
      .valid(valid),
      .h_cnt(h_cnt),
      .v_cnt(v_cnt)
    );
    
    /*wire flag;
    assign pass = (flag == 1'b1) ? 1'b1 : 1'b0;*/
    
    /*mem_addr_gen mem_addr_gen_inst(
    .clk(clk),
    .rst(rst),
    .hold(de_hold),
    .shift(shift_down),
    .rotate(rotate),
    .h_cnt(h_cnt),
    .v_cnt(v_cnt),
    .pixel_addr(pixel_addr),
    .flag(flag)
    );*/
parameter [14:0] state_0 [0:6399] = {
15'd0,15'd1,15'd2,15'd3,15'd4,15'd5,15'd6,15'd7,15'd8,15'd9,15'd10,15'd11,15'd12,15'd13,15'd14,15'd15,15'd16,15'd17,15'd18,15'd19,15'd20,15'd21,15'd22,15'd23,15'd24,15'd25,15'd26,15'd27,15'd28,15'd29,15'd30,15'd31,15'd32,15'd33,15'd34,15'd35,15'd36,15'd37,15'd38,15'd39,15'd40,15'd41,15'd42,15'd43,15'd44,15'd45,15'd46,15'd47,15'd48,15'd49,15'd50,15'd51,15'd52,15'd53,15'd54,15'd55,15'd56,15'd57,15'd58,15'd59,15'd60,15'd61,15'd62,15'd63,15'd64,15'd65,15'd66,15'd67,15'd68,15'd69,15'd70,15'd71,15'd72,15'd73,15'd74,15'd75,15'd76,15'd77,15'd78,15'd79,
15'd320,15'd321,15'd322,15'd323,15'd324,15'd325,15'd326,15'd327,15'd328,15'd329,15'd330,15'd331,15'd332,15'd333,15'd334,15'd335,15'd336,15'd337,15'd338,15'd339,15'd340,15'd341,15'd342,15'd343,15'd344,15'd345,15'd346,15'd347,15'd348,15'd349,15'd350,15'd351,15'd352,15'd353,15'd354,15'd355,15'd356,15'd357,15'd358,15'd359,15'd360,15'd361,15'd362,15'd363,15'd364,15'd365,15'd366,15'd367,15'd368,15'd369,15'd370,15'd371,15'd372,15'd373,15'd374,15'd375,15'd376,15'd377,15'd378,15'd379,15'd380,15'd381,15'd382,15'd383,15'd384,15'd385,15'd386,15'd387,15'd388,15'd389,15'd390,15'd391,15'd392,15'd393,15'd394,15'd395,15'd396,15'd397,15'd398,15'd399,
15'd640,15'd641,15'd642,15'd643,15'd644,15'd645,15'd646,15'd647,15'd648,15'd649,15'd650,15'd651,15'd652,15'd653,15'd654,15'd655,15'd656,15'd657,15'd658,15'd659,15'd660,15'd661,15'd662,15'd663,15'd664,15'd665,15'd666,15'd667,15'd668,15'd669,15'd670,15'd671,15'd672,15'd673,15'd674,15'd675,15'd676,15'd677,15'd678,15'd679,15'd680,15'd681,15'd682,15'd683,15'd684,15'd685,15'd686,15'd687,15'd688,15'd689,15'd690,15'd691,15'd692,15'd693,15'd694,15'd695,15'd696,15'd697,15'd698,15'd699,15'd700,15'd701,15'd702,15'd703,15'd704,15'd705,15'd706,15'd707,15'd708,15'd709,15'd710,15'd711,15'd712,15'd713,15'd714,15'd715,15'd716,15'd717,15'd718,15'd719,
15'd960,15'd961,15'd962,15'd963,15'd964,15'd965,15'd966,15'd967,15'd968,15'd969,15'd970,15'd971,15'd972,15'd973,15'd974,15'd975,15'd976,15'd977,15'd978,15'd979,15'd980,15'd981,15'd982,15'd983,15'd984,15'd985,15'd986,15'd987,15'd988,15'd989,15'd990,15'd991,15'd992,15'd993,15'd994,15'd995,15'd996,15'd997,15'd998,15'd999,15'd1000,15'd1001,15'd1002,15'd1003,15'd1004,15'd1005,15'd1006,15'd1007,15'd1008,15'd1009,15'd1010,15'd1011,15'd1012,15'd1013,15'd1014,15'd1015,15'd1016,15'd1017,15'd1018,15'd1019,15'd1020,15'd1021,15'd1022,15'd1023,15'd1024,15'd1025,15'd1026,15'd1027,15'd1028,15'd1029,15'd1030,15'd1031,15'd1032,15'd1033,15'd1034,15'd1035,15'd1036,15'd1037,15'd1038,15'd1039,
15'd1280,15'd1281,15'd1282,15'd1283,15'd1284,15'd1285,15'd1286,15'd1287,15'd1288,15'd1289,15'd1290,15'd1291,15'd1292,15'd1293,15'd1294,15'd1295,15'd1296,15'd1297,15'd1298,15'd1299,15'd1300,15'd1301,15'd1302,15'd1303,15'd1304,15'd1305,15'd1306,15'd1307,15'd1308,15'd1309,15'd1310,15'd1311,15'd1312,15'd1313,15'd1314,15'd1315,15'd1316,15'd1317,15'd1318,15'd1319,15'd1320,15'd1321,15'd1322,15'd1323,15'd1324,15'd1325,15'd1326,15'd1327,15'd1328,15'd1329,15'd1330,15'd1331,15'd1332,15'd1333,15'd1334,15'd1335,15'd1336,15'd1337,15'd1338,15'd1339,15'd1340,15'd1341,15'd1342,15'd1343,15'd1344,15'd1345,15'd1346,15'd1347,15'd1348,15'd1349,15'd1350,15'd1351,15'd1352,15'd1353,15'd1354,15'd1355,15'd1356,15'd1357,15'd1358,15'd1359,
15'd1600,15'd1601,15'd1602,15'd1603,15'd1604,15'd1605,15'd1606,15'd1607,15'd1608,15'd1609,15'd1610,15'd1611,15'd1612,15'd1613,15'd1614,15'd1615,15'd1616,15'd1617,15'd1618,15'd1619,15'd1620,15'd1621,15'd1622,15'd1623,15'd1624,15'd1625,15'd1626,15'd1627,15'd1628,15'd1629,15'd1630,15'd1631,15'd1632,15'd1633,15'd1634,15'd1635,15'd1636,15'd1637,15'd1638,15'd1639,15'd1640,15'd1641,15'd1642,15'd1643,15'd1644,15'd1645,15'd1646,15'd1647,15'd1648,15'd1649,15'd1650,15'd1651,15'd1652,15'd1653,15'd1654,15'd1655,15'd1656,15'd1657,15'd1658,15'd1659,15'd1660,15'd1661,15'd1662,15'd1663,15'd1664,15'd1665,15'd1666,15'd1667,15'd1668,15'd1669,15'd1670,15'd1671,15'd1672,15'd1673,15'd1674,15'd1675,15'd1676,15'd1677,15'd1678,15'd1679,
15'd1920,15'd1921,15'd1922,15'd1923,15'd1924,15'd1925,15'd1926,15'd1927,15'd1928,15'd1929,15'd1930,15'd1931,15'd1932,15'd1933,15'd1934,15'd1935,15'd1936,15'd1937,15'd1938,15'd1939,15'd1940,15'd1941,15'd1942,15'd1943,15'd1944,15'd1945,15'd1946,15'd1947,15'd1948,15'd1949,15'd1950,15'd1951,15'd1952,15'd1953,15'd1954,15'd1955,15'd1956,15'd1957,15'd1958,15'd1959,15'd1960,15'd1961,15'd1962,15'd1963,15'd1964,15'd1965,15'd1966,15'd1967,15'd1968,15'd1969,15'd1970,15'd1971,15'd1972,15'd1973,15'd1974,15'd1975,15'd1976,15'd1977,15'd1978,15'd1979,15'd1980,15'd1981,15'd1982,15'd1983,15'd1984,15'd1985,15'd1986,15'd1987,15'd1988,15'd1989,15'd1990,15'd1991,15'd1992,15'd1993,15'd1994,15'd1995,15'd1996,15'd1997,15'd1998,15'd1999,
15'd2240,15'd2241,15'd2242,15'd2243,15'd2244,15'd2245,15'd2246,15'd2247,15'd2248,15'd2249,15'd2250,15'd2251,15'd2252,15'd2253,15'd2254,15'd2255,15'd2256,15'd2257,15'd2258,15'd2259,15'd2260,15'd2261,15'd2262,15'd2263,15'd2264,15'd2265,15'd2266,15'd2267,15'd2268,15'd2269,15'd2270,15'd2271,15'd2272,15'd2273,15'd2274,15'd2275,15'd2276,15'd2277,15'd2278,15'd2279,15'd2280,15'd2281,15'd2282,15'd2283,15'd2284,15'd2285,15'd2286,15'd2287,15'd2288,15'd2289,15'd2290,15'd2291,15'd2292,15'd2293,15'd2294,15'd2295,15'd2296,15'd2297,15'd2298,15'd2299,15'd2300,15'd2301,15'd2302,15'd2303,15'd2304,15'd2305,15'd2306,15'd2307,15'd2308,15'd2309,15'd2310,15'd2311,15'd2312,15'd2313,15'd2314,15'd2315,15'd2316,15'd2317,15'd2318,15'd2319,
15'd2560,15'd2561,15'd2562,15'd2563,15'd2564,15'd2565,15'd2566,15'd2567,15'd2568,15'd2569,15'd2570,15'd2571,15'd2572,15'd2573,15'd2574,15'd2575,15'd2576,15'd2577,15'd2578,15'd2579,15'd2580,15'd2581,15'd2582,15'd2583,15'd2584,15'd2585,15'd2586,15'd2587,15'd2588,15'd2589,15'd2590,15'd2591,15'd2592,15'd2593,15'd2594,15'd2595,15'd2596,15'd2597,15'd2598,15'd2599,15'd2600,15'd2601,15'd2602,15'd2603,15'd2604,15'd2605,15'd2606,15'd2607,15'd2608,15'd2609,15'd2610,15'd2611,15'd2612,15'd2613,15'd2614,15'd2615,15'd2616,15'd2617,15'd2618,15'd2619,15'd2620,15'd2621,15'd2622,15'd2623,15'd2624,15'd2625,15'd2626,15'd2627,15'd2628,15'd2629,15'd2630,15'd2631,15'd2632,15'd2633,15'd2634,15'd2635,15'd2636,15'd2637,15'd2638,15'd2639,
15'd2880,15'd2881,15'd2882,15'd2883,15'd2884,15'd2885,15'd2886,15'd2887,15'd2888,15'd2889,15'd2890,15'd2891,15'd2892,15'd2893,15'd2894,15'd2895,15'd2896,15'd2897,15'd2898,15'd2899,15'd2900,15'd2901,15'd2902,15'd2903,15'd2904,15'd2905,15'd2906,15'd2907,15'd2908,15'd2909,15'd2910,15'd2911,15'd2912,15'd2913,15'd2914,15'd2915,15'd2916,15'd2917,15'd2918,15'd2919,15'd2920,15'd2921,15'd2922,15'd2923,15'd2924,15'd2925,15'd2926,15'd2927,15'd2928,15'd2929,15'd2930,15'd2931,15'd2932,15'd2933,15'd2934,15'd2935,15'd2936,15'd2937,15'd2938,15'd2939,15'd2940,15'd2941,15'd2942,15'd2943,15'd2944,15'd2945,15'd2946,15'd2947,15'd2948,15'd2949,15'd2950,15'd2951,15'd2952,15'd2953,15'd2954,15'd2955,15'd2956,15'd2957,15'd2958,15'd2959,
15'd3200,15'd3201,15'd3202,15'd3203,15'd3204,15'd3205,15'd3206,15'd3207,15'd3208,15'd3209,15'd3210,15'd3211,15'd3212,15'd3213,15'd3214,15'd3215,15'd3216,15'd3217,15'd3218,15'd3219,15'd3220,15'd3221,15'd3222,15'd3223,15'd3224,15'd3225,15'd3226,15'd3227,15'd3228,15'd3229,15'd3230,15'd3231,15'd3232,15'd3233,15'd3234,15'd3235,15'd3236,15'd3237,15'd3238,15'd3239,15'd3240,15'd3241,15'd3242,15'd3243,15'd3244,15'd3245,15'd3246,15'd3247,15'd3248,15'd3249,15'd3250,15'd3251,15'd3252,15'd3253,15'd3254,15'd3255,15'd3256,15'd3257,15'd3258,15'd3259,15'd3260,15'd3261,15'd3262,15'd3263,15'd3264,15'd3265,15'd3266,15'd3267,15'd3268,15'd3269,15'd3270,15'd3271,15'd3272,15'd3273,15'd3274,15'd3275,15'd3276,15'd3277,15'd3278,15'd3279,
15'd3520,15'd3521,15'd3522,15'd3523,15'd3524,15'd3525,15'd3526,15'd3527,15'd3528,15'd3529,15'd3530,15'd3531,15'd3532,15'd3533,15'd3534,15'd3535,15'd3536,15'd3537,15'd3538,15'd3539,15'd3540,15'd3541,15'd3542,15'd3543,15'd3544,15'd3545,15'd3546,15'd3547,15'd3548,15'd3549,15'd3550,15'd3551,15'd3552,15'd3553,15'd3554,15'd3555,15'd3556,15'd3557,15'd3558,15'd3559,15'd3560,15'd3561,15'd3562,15'd3563,15'd3564,15'd3565,15'd3566,15'd3567,15'd3568,15'd3569,15'd3570,15'd3571,15'd3572,15'd3573,15'd3574,15'd3575,15'd3576,15'd3577,15'd3578,15'd3579,15'd3580,15'd3581,15'd3582,15'd3583,15'd3584,15'd3585,15'd3586,15'd3587,15'd3588,15'd3589,15'd3590,15'd3591,15'd3592,15'd3593,15'd3594,15'd3595,15'd3596,15'd3597,15'd3598,15'd3599,
15'd3840,15'd3841,15'd3842,15'd3843,15'd3844,15'd3845,15'd3846,15'd3847,15'd3848,15'd3849,15'd3850,15'd3851,15'd3852,15'd3853,15'd3854,15'd3855,15'd3856,15'd3857,15'd3858,15'd3859,15'd3860,15'd3861,15'd3862,15'd3863,15'd3864,15'd3865,15'd3866,15'd3867,15'd3868,15'd3869,15'd3870,15'd3871,15'd3872,15'd3873,15'd3874,15'd3875,15'd3876,15'd3877,15'd3878,15'd3879,15'd3880,15'd3881,15'd3882,15'd3883,15'd3884,15'd3885,15'd3886,15'd3887,15'd3888,15'd3889,15'd3890,15'd3891,15'd3892,15'd3893,15'd3894,15'd3895,15'd3896,15'd3897,15'd3898,15'd3899,15'd3900,15'd3901,15'd3902,15'd3903,15'd3904,15'd3905,15'd3906,15'd3907,15'd3908,15'd3909,15'd3910,15'd3911,15'd3912,15'd3913,15'd3914,15'd3915,15'd3916,15'd3917,15'd3918,15'd3919,
15'd4160,15'd4161,15'd4162,15'd4163,15'd4164,15'd4165,15'd4166,15'd4167,15'd4168,15'd4169,15'd4170,15'd4171,15'd4172,15'd4173,15'd4174,15'd4175,15'd4176,15'd4177,15'd4178,15'd4179,15'd4180,15'd4181,15'd4182,15'd4183,15'd4184,15'd4185,15'd4186,15'd4187,15'd4188,15'd4189,15'd4190,15'd4191,15'd4192,15'd4193,15'd4194,15'd4195,15'd4196,15'd4197,15'd4198,15'd4199,15'd4200,15'd4201,15'd4202,15'd4203,15'd4204,15'd4205,15'd4206,15'd4207,15'd4208,15'd4209,15'd4210,15'd4211,15'd4212,15'd4213,15'd4214,15'd4215,15'd4216,15'd4217,15'd4218,15'd4219,15'd4220,15'd4221,15'd4222,15'd4223,15'd4224,15'd4225,15'd4226,15'd4227,15'd4228,15'd4229,15'd4230,15'd4231,15'd4232,15'd4233,15'd4234,15'd4235,15'd4236,15'd4237,15'd4238,15'd4239,
15'd4480,15'd4481,15'd4482,15'd4483,15'd4484,15'd4485,15'd4486,15'd4487,15'd4488,15'd4489,15'd4490,15'd4491,15'd4492,15'd4493,15'd4494,15'd4495,15'd4496,15'd4497,15'd4498,15'd4499,15'd4500,15'd4501,15'd4502,15'd4503,15'd4504,15'd4505,15'd4506,15'd4507,15'd4508,15'd4509,15'd4510,15'd4511,15'd4512,15'd4513,15'd4514,15'd4515,15'd4516,15'd4517,15'd4518,15'd4519,15'd4520,15'd4521,15'd4522,15'd4523,15'd4524,15'd4525,15'd4526,15'd4527,15'd4528,15'd4529,15'd4530,15'd4531,15'd4532,15'd4533,15'd4534,15'd4535,15'd4536,15'd4537,15'd4538,15'd4539,15'd4540,15'd4541,15'd4542,15'd4543,15'd4544,15'd4545,15'd4546,15'd4547,15'd4548,15'd4549,15'd4550,15'd4551,15'd4552,15'd4553,15'd4554,15'd4555,15'd4556,15'd4557,15'd4558,15'd4559,
15'd4800,15'd4801,15'd4802,15'd4803,15'd4804,15'd4805,15'd4806,15'd4807,15'd4808,15'd4809,15'd4810,15'd4811,15'd4812,15'd4813,15'd4814,15'd4815,15'd4816,15'd4817,15'd4818,15'd4819,15'd4820,15'd4821,15'd4822,15'd4823,15'd4824,15'd4825,15'd4826,15'd4827,15'd4828,15'd4829,15'd4830,15'd4831,15'd4832,15'd4833,15'd4834,15'd4835,15'd4836,15'd4837,15'd4838,15'd4839,15'd4840,15'd4841,15'd4842,15'd4843,15'd4844,15'd4845,15'd4846,15'd4847,15'd4848,15'd4849,15'd4850,15'd4851,15'd4852,15'd4853,15'd4854,15'd4855,15'd4856,15'd4857,15'd4858,15'd4859,15'd4860,15'd4861,15'd4862,15'd4863,15'd4864,15'd4865,15'd4866,15'd4867,15'd4868,15'd4869,15'd4870,15'd4871,15'd4872,15'd4873,15'd4874,15'd4875,15'd4876,15'd4877,15'd4878,15'd4879,
15'd5120,15'd5121,15'd5122,15'd5123,15'd5124,15'd5125,15'd5126,15'd5127,15'd5128,15'd5129,15'd5130,15'd5131,15'd5132,15'd5133,15'd5134,15'd5135,15'd5136,15'd5137,15'd5138,15'd5139,15'd5140,15'd5141,15'd5142,15'd5143,15'd5144,15'd5145,15'd5146,15'd5147,15'd5148,15'd5149,15'd5150,15'd5151,15'd5152,15'd5153,15'd5154,15'd5155,15'd5156,15'd5157,15'd5158,15'd5159,15'd5160,15'd5161,15'd5162,15'd5163,15'd5164,15'd5165,15'd5166,15'd5167,15'd5168,15'd5169,15'd5170,15'd5171,15'd5172,15'd5173,15'd5174,15'd5175,15'd5176,15'd5177,15'd5178,15'd5179,15'd5180,15'd5181,15'd5182,15'd5183,15'd5184,15'd5185,15'd5186,15'd5187,15'd5188,15'd5189,15'd5190,15'd5191,15'd5192,15'd5193,15'd5194,15'd5195,15'd5196,15'd5197,15'd5198,15'd5199,
15'd5440,15'd5441,15'd5442,15'd5443,15'd5444,15'd5445,15'd5446,15'd5447,15'd5448,15'd5449,15'd5450,15'd5451,15'd5452,15'd5453,15'd5454,15'd5455,15'd5456,15'd5457,15'd5458,15'd5459,15'd5460,15'd5461,15'd5462,15'd5463,15'd5464,15'd5465,15'd5466,15'd5467,15'd5468,15'd5469,15'd5470,15'd5471,15'd5472,15'd5473,15'd5474,15'd5475,15'd5476,15'd5477,15'd5478,15'd5479,15'd5480,15'd5481,15'd5482,15'd5483,15'd5484,15'd5485,15'd5486,15'd5487,15'd5488,15'd5489,15'd5490,15'd5491,15'd5492,15'd5493,15'd5494,15'd5495,15'd5496,15'd5497,15'd5498,15'd5499,15'd5500,15'd5501,15'd5502,15'd5503,15'd5504,15'd5505,15'd5506,15'd5507,15'd5508,15'd5509,15'd5510,15'd5511,15'd5512,15'd5513,15'd5514,15'd5515,15'd5516,15'd5517,15'd5518,15'd5519,
15'd5760,15'd5761,15'd5762,15'd5763,15'd5764,15'd5765,15'd5766,15'd5767,15'd5768,15'd5769,15'd5770,15'd5771,15'd5772,15'd5773,15'd5774,15'd5775,15'd5776,15'd5777,15'd5778,15'd5779,15'd5780,15'd5781,15'd5782,15'd5783,15'd5784,15'd5785,15'd5786,15'd5787,15'd5788,15'd5789,15'd5790,15'd5791,15'd5792,15'd5793,15'd5794,15'd5795,15'd5796,15'd5797,15'd5798,15'd5799,15'd5800,15'd5801,15'd5802,15'd5803,15'd5804,15'd5805,15'd5806,15'd5807,15'd5808,15'd5809,15'd5810,15'd5811,15'd5812,15'd5813,15'd5814,15'd5815,15'd5816,15'd5817,15'd5818,15'd5819,15'd5820,15'd5821,15'd5822,15'd5823,15'd5824,15'd5825,15'd5826,15'd5827,15'd5828,15'd5829,15'd5830,15'd5831,15'd5832,15'd5833,15'd5834,15'd5835,15'd5836,15'd5837,15'd5838,15'd5839,
15'd6080,15'd6081,15'd6082,15'd6083,15'd6084,15'd6085,15'd6086,15'd6087,15'd6088,15'd6089,15'd6090,15'd6091,15'd6092,15'd6093,15'd6094,15'd6095,15'd6096,15'd6097,15'd6098,15'd6099,15'd6100,15'd6101,15'd6102,15'd6103,15'd6104,15'd6105,15'd6106,15'd6107,15'd6108,15'd6109,15'd6110,15'd6111,15'd6112,15'd6113,15'd6114,15'd6115,15'd6116,15'd6117,15'd6118,15'd6119,15'd6120,15'd6121,15'd6122,15'd6123,15'd6124,15'd6125,15'd6126,15'd6127,15'd6128,15'd6129,15'd6130,15'd6131,15'd6132,15'd6133,15'd6134,15'd6135,15'd6136,15'd6137,15'd6138,15'd6139,15'd6140,15'd6141,15'd6142,15'd6143,15'd6144,15'd6145,15'd6146,15'd6147,15'd6148,15'd6149,15'd6150,15'd6151,15'd6152,15'd6153,15'd6154,15'd6155,15'd6156,15'd6157,15'd6158,15'd6159,
15'd6400,15'd6401,15'd6402,15'd6403,15'd6404,15'd6405,15'd6406,15'd6407,15'd6408,15'd6409,15'd6410,15'd6411,15'd6412,15'd6413,15'd6414,15'd6415,15'd6416,15'd6417,15'd6418,15'd6419,15'd6420,15'd6421,15'd6422,15'd6423,15'd6424,15'd6425,15'd6426,15'd6427,15'd6428,15'd6429,15'd6430,15'd6431,15'd6432,15'd6433,15'd6434,15'd6435,15'd6436,15'd6437,15'd6438,15'd6439,15'd6440,15'd6441,15'd6442,15'd6443,15'd6444,15'd6445,15'd6446,15'd6447,15'd6448,15'd6449,15'd6450,15'd6451,15'd6452,15'd6453,15'd6454,15'd6455,15'd6456,15'd6457,15'd6458,15'd6459,15'd6460,15'd6461,15'd6462,15'd6463,15'd6464,15'd6465,15'd6466,15'd6467,15'd6468,15'd6469,15'd6470,15'd6471,15'd6472,15'd6473,15'd6474,15'd6475,15'd6476,15'd6477,15'd6478,15'd6479,
15'd6720,15'd6721,15'd6722,15'd6723,15'd6724,15'd6725,15'd6726,15'd6727,15'd6728,15'd6729,15'd6730,15'd6731,15'd6732,15'd6733,15'd6734,15'd6735,15'd6736,15'd6737,15'd6738,15'd6739,15'd6740,15'd6741,15'd6742,15'd6743,15'd6744,15'd6745,15'd6746,15'd6747,15'd6748,15'd6749,15'd6750,15'd6751,15'd6752,15'd6753,15'd6754,15'd6755,15'd6756,15'd6757,15'd6758,15'd6759,15'd6760,15'd6761,15'd6762,15'd6763,15'd6764,15'd6765,15'd6766,15'd6767,15'd6768,15'd6769,15'd6770,15'd6771,15'd6772,15'd6773,15'd6774,15'd6775,15'd6776,15'd6777,15'd6778,15'd6779,15'd6780,15'd6781,15'd6782,15'd6783,15'd6784,15'd6785,15'd6786,15'd6787,15'd6788,15'd6789,15'd6790,15'd6791,15'd6792,15'd6793,15'd6794,15'd6795,15'd6796,15'd6797,15'd6798,15'd6799,
15'd7040,15'd7041,15'd7042,15'd7043,15'd7044,15'd7045,15'd7046,15'd7047,15'd7048,15'd7049,15'd7050,15'd7051,15'd7052,15'd7053,15'd7054,15'd7055,15'd7056,15'd7057,15'd7058,15'd7059,15'd7060,15'd7061,15'd7062,15'd7063,15'd7064,15'd7065,15'd7066,15'd7067,15'd7068,15'd7069,15'd7070,15'd7071,15'd7072,15'd7073,15'd7074,15'd7075,15'd7076,15'd7077,15'd7078,15'd7079,15'd7080,15'd7081,15'd7082,15'd7083,15'd7084,15'd7085,15'd7086,15'd7087,15'd7088,15'd7089,15'd7090,15'd7091,15'd7092,15'd7093,15'd7094,15'd7095,15'd7096,15'd7097,15'd7098,15'd7099,15'd7100,15'd7101,15'd7102,15'd7103,15'd7104,15'd7105,15'd7106,15'd7107,15'd7108,15'd7109,15'd7110,15'd7111,15'd7112,15'd7113,15'd7114,15'd7115,15'd7116,15'd7117,15'd7118,15'd7119,
15'd7360,15'd7361,15'd7362,15'd7363,15'd7364,15'd7365,15'd7366,15'd7367,15'd7368,15'd7369,15'd7370,15'd7371,15'd7372,15'd7373,15'd7374,15'd7375,15'd7376,15'd7377,15'd7378,15'd7379,15'd7380,15'd7381,15'd7382,15'd7383,15'd7384,15'd7385,15'd7386,15'd7387,15'd7388,15'd7389,15'd7390,15'd7391,15'd7392,15'd7393,15'd7394,15'd7395,15'd7396,15'd7397,15'd7398,15'd7399,15'd7400,15'd7401,15'd7402,15'd7403,15'd7404,15'd7405,15'd7406,15'd7407,15'd7408,15'd7409,15'd7410,15'd7411,15'd7412,15'd7413,15'd7414,15'd7415,15'd7416,15'd7417,15'd7418,15'd7419,15'd7420,15'd7421,15'd7422,15'd7423,15'd7424,15'd7425,15'd7426,15'd7427,15'd7428,15'd7429,15'd7430,15'd7431,15'd7432,15'd7433,15'd7434,15'd7435,15'd7436,15'd7437,15'd7438,15'd7439,
15'd7680,15'd7681,15'd7682,15'd7683,15'd7684,15'd7685,15'd7686,15'd7687,15'd7688,15'd7689,15'd7690,15'd7691,15'd7692,15'd7693,15'd7694,15'd7695,15'd7696,15'd7697,15'd7698,15'd7699,15'd7700,15'd7701,15'd7702,15'd7703,15'd7704,15'd7705,15'd7706,15'd7707,15'd7708,15'd7709,15'd7710,15'd7711,15'd7712,15'd7713,15'd7714,15'd7715,15'd7716,15'd7717,15'd7718,15'd7719,15'd7720,15'd7721,15'd7722,15'd7723,15'd7724,15'd7725,15'd7726,15'd7727,15'd7728,15'd7729,15'd7730,15'd7731,15'd7732,15'd7733,15'd7734,15'd7735,15'd7736,15'd7737,15'd7738,15'd7739,15'd7740,15'd7741,15'd7742,15'd7743,15'd7744,15'd7745,15'd7746,15'd7747,15'd7748,15'd7749,15'd7750,15'd7751,15'd7752,15'd7753,15'd7754,15'd7755,15'd7756,15'd7757,15'd7758,15'd7759,
15'd8000,15'd8001,15'd8002,15'd8003,15'd8004,15'd8005,15'd8006,15'd8007,15'd8008,15'd8009,15'd8010,15'd8011,15'd8012,15'd8013,15'd8014,15'd8015,15'd8016,15'd8017,15'd8018,15'd8019,15'd8020,15'd8021,15'd8022,15'd8023,15'd8024,15'd8025,15'd8026,15'd8027,15'd8028,15'd8029,15'd8030,15'd8031,15'd8032,15'd8033,15'd8034,15'd8035,15'd8036,15'd8037,15'd8038,15'd8039,15'd8040,15'd8041,15'd8042,15'd8043,15'd8044,15'd8045,15'd8046,15'd8047,15'd8048,15'd8049,15'd8050,15'd8051,15'd8052,15'd8053,15'd8054,15'd8055,15'd8056,15'd8057,15'd8058,15'd8059,15'd8060,15'd8061,15'd8062,15'd8063,15'd8064,15'd8065,15'd8066,15'd8067,15'd8068,15'd8069,15'd8070,15'd8071,15'd8072,15'd8073,15'd8074,15'd8075,15'd8076,15'd8077,15'd8078,15'd8079,
15'd8320,15'd8321,15'd8322,15'd8323,15'd8324,15'd8325,15'd8326,15'd8327,15'd8328,15'd8329,15'd8330,15'd8331,15'd8332,15'd8333,15'd8334,15'd8335,15'd8336,15'd8337,15'd8338,15'd8339,15'd8340,15'd8341,15'd8342,15'd8343,15'd8344,15'd8345,15'd8346,15'd8347,15'd8348,15'd8349,15'd8350,15'd8351,15'd8352,15'd8353,15'd8354,15'd8355,15'd8356,15'd8357,15'd8358,15'd8359,15'd8360,15'd8361,15'd8362,15'd8363,15'd8364,15'd8365,15'd8366,15'd8367,15'd8368,15'd8369,15'd8370,15'd8371,15'd8372,15'd8373,15'd8374,15'd8375,15'd8376,15'd8377,15'd8378,15'd8379,15'd8380,15'd8381,15'd8382,15'd8383,15'd8384,15'd8385,15'd8386,15'd8387,15'd8388,15'd8389,15'd8390,15'd8391,15'd8392,15'd8393,15'd8394,15'd8395,15'd8396,15'd8397,15'd8398,15'd8399,
15'd8640,15'd8641,15'd8642,15'd8643,15'd8644,15'd8645,15'd8646,15'd8647,15'd8648,15'd8649,15'd8650,15'd8651,15'd8652,15'd8653,15'd8654,15'd8655,15'd8656,15'd8657,15'd8658,15'd8659,15'd8660,15'd8661,15'd8662,15'd8663,15'd8664,15'd8665,15'd8666,15'd8667,15'd8668,15'd8669,15'd8670,15'd8671,15'd8672,15'd8673,15'd8674,15'd8675,15'd8676,15'd8677,15'd8678,15'd8679,15'd8680,15'd8681,15'd8682,15'd8683,15'd8684,15'd8685,15'd8686,15'd8687,15'd8688,15'd8689,15'd8690,15'd8691,15'd8692,15'd8693,15'd8694,15'd8695,15'd8696,15'd8697,15'd8698,15'd8699,15'd8700,15'd8701,15'd8702,15'd8703,15'd8704,15'd8705,15'd8706,15'd8707,15'd8708,15'd8709,15'd8710,15'd8711,15'd8712,15'd8713,15'd8714,15'd8715,15'd8716,15'd8717,15'd8718,15'd8719,
15'd8960,15'd8961,15'd8962,15'd8963,15'd8964,15'd8965,15'd8966,15'd8967,15'd8968,15'd8969,15'd8970,15'd8971,15'd8972,15'd8973,15'd8974,15'd8975,15'd8976,15'd8977,15'd8978,15'd8979,15'd8980,15'd8981,15'd8982,15'd8983,15'd8984,15'd8985,15'd8986,15'd8987,15'd8988,15'd8989,15'd8990,15'd8991,15'd8992,15'd8993,15'd8994,15'd8995,15'd8996,15'd8997,15'd8998,15'd8999,15'd9000,15'd9001,15'd9002,15'd9003,15'd9004,15'd9005,15'd9006,15'd9007,15'd9008,15'd9009,15'd9010,15'd9011,15'd9012,15'd9013,15'd9014,15'd9015,15'd9016,15'd9017,15'd9018,15'd9019,15'd9020,15'd9021,15'd9022,15'd9023,15'd9024,15'd9025,15'd9026,15'd9027,15'd9028,15'd9029,15'd9030,15'd9031,15'd9032,15'd9033,15'd9034,15'd9035,15'd9036,15'd9037,15'd9038,15'd9039,
15'd9280,15'd9281,15'd9282,15'd9283,15'd9284,15'd9285,15'd9286,15'd9287,15'd9288,15'd9289,15'd9290,15'd9291,15'd9292,15'd9293,15'd9294,15'd9295,15'd9296,15'd9297,15'd9298,15'd9299,15'd9300,15'd9301,15'd9302,15'd9303,15'd9304,15'd9305,15'd9306,15'd9307,15'd9308,15'd9309,15'd9310,15'd9311,15'd9312,15'd9313,15'd9314,15'd9315,15'd9316,15'd9317,15'd9318,15'd9319,15'd9320,15'd9321,15'd9322,15'd9323,15'd9324,15'd9325,15'd9326,15'd9327,15'd9328,15'd9329,15'd9330,15'd9331,15'd9332,15'd9333,15'd9334,15'd9335,15'd9336,15'd9337,15'd9338,15'd9339,15'd9340,15'd9341,15'd9342,15'd9343,15'd9344,15'd9345,15'd9346,15'd9347,15'd9348,15'd9349,15'd9350,15'd9351,15'd9352,15'd9353,15'd9354,15'd9355,15'd9356,15'd9357,15'd9358,15'd9359,
15'd9600,15'd9601,15'd9602,15'd9603,15'd9604,15'd9605,15'd9606,15'd9607,15'd9608,15'd9609,15'd9610,15'd9611,15'd9612,15'd9613,15'd9614,15'd9615,15'd9616,15'd9617,15'd9618,15'd9619,15'd9620,15'd9621,15'd9622,15'd9623,15'd9624,15'd9625,15'd9626,15'd9627,15'd9628,15'd9629,15'd9630,15'd9631,15'd9632,15'd9633,15'd9634,15'd9635,15'd9636,15'd9637,15'd9638,15'd9639,15'd9640,15'd9641,15'd9642,15'd9643,15'd9644,15'd9645,15'd9646,15'd9647,15'd9648,15'd9649,15'd9650,15'd9651,15'd9652,15'd9653,15'd9654,15'd9655,15'd9656,15'd9657,15'd9658,15'd9659,15'd9660,15'd9661,15'd9662,15'd9663,15'd9664,15'd9665,15'd9666,15'd9667,15'd9668,15'd9669,15'd9670,15'd9671,15'd9672,15'd9673,15'd9674,15'd9675,15'd9676,15'd9677,15'd9678,15'd9679,
15'd9920,15'd9921,15'd9922,15'd9923,15'd9924,15'd9925,15'd9926,15'd9927,15'd9928,15'd9929,15'd9930,15'd9931,15'd9932,15'd9933,15'd9934,15'd9935,15'd9936,15'd9937,15'd9938,15'd9939,15'd9940,15'd9941,15'd9942,15'd9943,15'd9944,15'd9945,15'd9946,15'd9947,15'd9948,15'd9949,15'd9950,15'd9951,15'd9952,15'd9953,15'd9954,15'd9955,15'd9956,15'd9957,15'd9958,15'd9959,15'd9960,15'd9961,15'd9962,15'd9963,15'd9964,15'd9965,15'd9966,15'd9967,15'd9968,15'd9969,15'd9970,15'd9971,15'd9972,15'd9973,15'd9974,15'd9975,15'd9976,15'd9977,15'd9978,15'd9979,15'd9980,15'd9981,15'd9982,15'd9983,15'd9984,15'd9985,15'd9986,15'd9987,15'd9988,15'd9989,15'd9990,15'd9991,15'd9992,15'd9993,15'd9994,15'd9995,15'd9996,15'd9997,15'd9998,15'd9999,
15'd10240,15'd10241,15'd10242,15'd10243,15'd10244,15'd10245,15'd10246,15'd10247,15'd10248,15'd10249,15'd10250,15'd10251,15'd10252,15'd10253,15'd10254,15'd10255,15'd10256,15'd10257,15'd10258,15'd10259,15'd10260,15'd10261,15'd10262,15'd10263,15'd10264,15'd10265,15'd10266,15'd10267,15'd10268,15'd10269,15'd10270,15'd10271,15'd10272,15'd10273,15'd10274,15'd10275,15'd10276,15'd10277,15'd10278,15'd10279,15'd10280,15'd10281,15'd10282,15'd10283,15'd10284,15'd10285,15'd10286,15'd10287,15'd10288,15'd10289,15'd10290,15'd10291,15'd10292,15'd10293,15'd10294,15'd10295,15'd10296,15'd10297,15'd10298,15'd10299,15'd10300,15'd10301,15'd10302,15'd10303,15'd10304,15'd10305,15'd10306,15'd10307,15'd10308,15'd10309,15'd10310,15'd10311,15'd10312,15'd10313,15'd10314,15'd10315,15'd10316,15'd10317,15'd10318,15'd10319,
15'd10560,15'd10561,15'd10562,15'd10563,15'd10564,15'd10565,15'd10566,15'd10567,15'd10568,15'd10569,15'd10570,15'd10571,15'd10572,15'd10573,15'd10574,15'd10575,15'd10576,15'd10577,15'd10578,15'd10579,15'd10580,15'd10581,15'd10582,15'd10583,15'd10584,15'd10585,15'd10586,15'd10587,15'd10588,15'd10589,15'd10590,15'd10591,15'd10592,15'd10593,15'd10594,15'd10595,15'd10596,15'd10597,15'd10598,15'd10599,15'd10600,15'd10601,15'd10602,15'd10603,15'd10604,15'd10605,15'd10606,15'd10607,15'd10608,15'd10609,15'd10610,15'd10611,15'd10612,15'd10613,15'd10614,15'd10615,15'd10616,15'd10617,15'd10618,15'd10619,15'd10620,15'd10621,15'd10622,15'd10623,15'd10624,15'd10625,15'd10626,15'd10627,15'd10628,15'd10629,15'd10630,15'd10631,15'd10632,15'd10633,15'd10634,15'd10635,15'd10636,15'd10637,15'd10638,15'd10639,
15'd10880,15'd10881,15'd10882,15'd10883,15'd10884,15'd10885,15'd10886,15'd10887,15'd10888,15'd10889,15'd10890,15'd10891,15'd10892,15'd10893,15'd10894,15'd10895,15'd10896,15'd10897,15'd10898,15'd10899,15'd10900,15'd10901,15'd10902,15'd10903,15'd10904,15'd10905,15'd10906,15'd10907,15'd10908,15'd10909,15'd10910,15'd10911,15'd10912,15'd10913,15'd10914,15'd10915,15'd10916,15'd10917,15'd10918,15'd10919,15'd10920,15'd10921,15'd10922,15'd10923,15'd10924,15'd10925,15'd10926,15'd10927,15'd10928,15'd10929,15'd10930,15'd10931,15'd10932,15'd10933,15'd10934,15'd10935,15'd10936,15'd10937,15'd10938,15'd10939,15'd10940,15'd10941,15'd10942,15'd10943,15'd10944,15'd10945,15'd10946,15'd10947,15'd10948,15'd10949,15'd10950,15'd10951,15'd10952,15'd10953,15'd10954,15'd10955,15'd10956,15'd10957,15'd10958,15'd10959,
15'd11200,15'd11201,15'd11202,15'd11203,15'd11204,15'd11205,15'd11206,15'd11207,15'd11208,15'd11209,15'd11210,15'd11211,15'd11212,15'd11213,15'd11214,15'd11215,15'd11216,15'd11217,15'd11218,15'd11219,15'd11220,15'd11221,15'd11222,15'd11223,15'd11224,15'd11225,15'd11226,15'd11227,15'd11228,15'd11229,15'd11230,15'd11231,15'd11232,15'd11233,15'd11234,15'd11235,15'd11236,15'd11237,15'd11238,15'd11239,15'd11240,15'd11241,15'd11242,15'd11243,15'd11244,15'd11245,15'd11246,15'd11247,15'd11248,15'd11249,15'd11250,15'd11251,15'd11252,15'd11253,15'd11254,15'd11255,15'd11256,15'd11257,15'd11258,15'd11259,15'd11260,15'd11261,15'd11262,15'd11263,15'd11264,15'd11265,15'd11266,15'd11267,15'd11268,15'd11269,15'd11270,15'd11271,15'd11272,15'd11273,15'd11274,15'd11275,15'd11276,15'd11277,15'd11278,15'd11279,
15'd11520,15'd11521,15'd11522,15'd11523,15'd11524,15'd11525,15'd11526,15'd11527,15'd11528,15'd11529,15'd11530,15'd11531,15'd11532,15'd11533,15'd11534,15'd11535,15'd11536,15'd11537,15'd11538,15'd11539,15'd11540,15'd11541,15'd11542,15'd11543,15'd11544,15'd11545,15'd11546,15'd11547,15'd11548,15'd11549,15'd11550,15'd11551,15'd11552,15'd11553,15'd11554,15'd11555,15'd11556,15'd11557,15'd11558,15'd11559,15'd11560,15'd11561,15'd11562,15'd11563,15'd11564,15'd11565,15'd11566,15'd11567,15'd11568,15'd11569,15'd11570,15'd11571,15'd11572,15'd11573,15'd11574,15'd11575,15'd11576,15'd11577,15'd11578,15'd11579,15'd11580,15'd11581,15'd11582,15'd11583,15'd11584,15'd11585,15'd11586,15'd11587,15'd11588,15'd11589,15'd11590,15'd11591,15'd11592,15'd11593,15'd11594,15'd11595,15'd11596,15'd11597,15'd11598,15'd11599,
15'd11840,15'd11841,15'd11842,15'd11843,15'd11844,15'd11845,15'd11846,15'd11847,15'd11848,15'd11849,15'd11850,15'd11851,15'd11852,15'd11853,15'd11854,15'd11855,15'd11856,15'd11857,15'd11858,15'd11859,15'd11860,15'd11861,15'd11862,15'd11863,15'd11864,15'd11865,15'd11866,15'd11867,15'd11868,15'd11869,15'd11870,15'd11871,15'd11872,15'd11873,15'd11874,15'd11875,15'd11876,15'd11877,15'd11878,15'd11879,15'd11880,15'd11881,15'd11882,15'd11883,15'd11884,15'd11885,15'd11886,15'd11887,15'd11888,15'd11889,15'd11890,15'd11891,15'd11892,15'd11893,15'd11894,15'd11895,15'd11896,15'd11897,15'd11898,15'd11899,15'd11900,15'd11901,15'd11902,15'd11903,15'd11904,15'd11905,15'd11906,15'd11907,15'd11908,15'd11909,15'd11910,15'd11911,15'd11912,15'd11913,15'd11914,15'd11915,15'd11916,15'd11917,15'd11918,15'd11919,
15'd12160,15'd12161,15'd12162,15'd12163,15'd12164,15'd12165,15'd12166,15'd12167,15'd12168,15'd12169,15'd12170,15'd12171,15'd12172,15'd12173,15'd12174,15'd12175,15'd12176,15'd12177,15'd12178,15'd12179,15'd12180,15'd12181,15'd12182,15'd12183,15'd12184,15'd12185,15'd12186,15'd12187,15'd12188,15'd12189,15'd12190,15'd12191,15'd12192,15'd12193,15'd12194,15'd12195,15'd12196,15'd12197,15'd12198,15'd12199,15'd12200,15'd12201,15'd12202,15'd12203,15'd12204,15'd12205,15'd12206,15'd12207,15'd12208,15'd12209,15'd12210,15'd12211,15'd12212,15'd12213,15'd12214,15'd12215,15'd12216,15'd12217,15'd12218,15'd12219,15'd12220,15'd12221,15'd12222,15'd12223,15'd12224,15'd12225,15'd12226,15'd12227,15'd12228,15'd12229,15'd12230,15'd12231,15'd12232,15'd12233,15'd12234,15'd12235,15'd12236,15'd12237,15'd12238,15'd12239,
15'd12480,15'd12481,15'd12482,15'd12483,15'd12484,15'd12485,15'd12486,15'd12487,15'd12488,15'd12489,15'd12490,15'd12491,15'd12492,15'd12493,15'd12494,15'd12495,15'd12496,15'd12497,15'd12498,15'd12499,15'd12500,15'd12501,15'd12502,15'd12503,15'd12504,15'd12505,15'd12506,15'd12507,15'd12508,15'd12509,15'd12510,15'd12511,15'd12512,15'd12513,15'd12514,15'd12515,15'd12516,15'd12517,15'd12518,15'd12519,15'd12520,15'd12521,15'd12522,15'd12523,15'd12524,15'd12525,15'd12526,15'd12527,15'd12528,15'd12529,15'd12530,15'd12531,15'd12532,15'd12533,15'd12534,15'd12535,15'd12536,15'd12537,15'd12538,15'd12539,15'd12540,15'd12541,15'd12542,15'd12543,15'd12544,15'd12545,15'd12546,15'd12547,15'd12548,15'd12549,15'd12550,15'd12551,15'd12552,15'd12553,15'd12554,15'd12555,15'd12556,15'd12557,15'd12558,15'd12559,
15'd12800,15'd12801,15'd12802,15'd12803,15'd12804,15'd12805,15'd12806,15'd12807,15'd12808,15'd12809,15'd12810,15'd12811,15'd12812,15'd12813,15'd12814,15'd12815,15'd12816,15'd12817,15'd12818,15'd12819,15'd12820,15'd12821,15'd12822,15'd12823,15'd12824,15'd12825,15'd12826,15'd12827,15'd12828,15'd12829,15'd12830,15'd12831,15'd12832,15'd12833,15'd12834,15'd12835,15'd12836,15'd12837,15'd12838,15'd12839,15'd12840,15'd12841,15'd12842,15'd12843,15'd12844,15'd12845,15'd12846,15'd12847,15'd12848,15'd12849,15'd12850,15'd12851,15'd12852,15'd12853,15'd12854,15'd12855,15'd12856,15'd12857,15'd12858,15'd12859,15'd12860,15'd12861,15'd12862,15'd12863,15'd12864,15'd12865,15'd12866,15'd12867,15'd12868,15'd12869,15'd12870,15'd12871,15'd12872,15'd12873,15'd12874,15'd12875,15'd12876,15'd12877,15'd12878,15'd12879,
15'd13120,15'd13121,15'd13122,15'd13123,15'd13124,15'd13125,15'd13126,15'd13127,15'd13128,15'd13129,15'd13130,15'd13131,15'd13132,15'd13133,15'd13134,15'd13135,15'd13136,15'd13137,15'd13138,15'd13139,15'd13140,15'd13141,15'd13142,15'd13143,15'd13144,15'd13145,15'd13146,15'd13147,15'd13148,15'd13149,15'd13150,15'd13151,15'd13152,15'd13153,15'd13154,15'd13155,15'd13156,15'd13157,15'd13158,15'd13159,15'd13160,15'd13161,15'd13162,15'd13163,15'd13164,15'd13165,15'd13166,15'd13167,15'd13168,15'd13169,15'd13170,15'd13171,15'd13172,15'd13173,15'd13174,15'd13175,15'd13176,15'd13177,15'd13178,15'd13179,15'd13180,15'd13181,15'd13182,15'd13183,15'd13184,15'd13185,15'd13186,15'd13187,15'd13188,15'd13189,15'd13190,15'd13191,15'd13192,15'd13193,15'd13194,15'd13195,15'd13196,15'd13197,15'd13198,15'd13199,
15'd13440,15'd13441,15'd13442,15'd13443,15'd13444,15'd13445,15'd13446,15'd13447,15'd13448,15'd13449,15'd13450,15'd13451,15'd13452,15'd13453,15'd13454,15'd13455,15'd13456,15'd13457,15'd13458,15'd13459,15'd13460,15'd13461,15'd13462,15'd13463,15'd13464,15'd13465,15'd13466,15'd13467,15'd13468,15'd13469,15'd13470,15'd13471,15'd13472,15'd13473,15'd13474,15'd13475,15'd13476,15'd13477,15'd13478,15'd13479,15'd13480,15'd13481,15'd13482,15'd13483,15'd13484,15'd13485,15'd13486,15'd13487,15'd13488,15'd13489,15'd13490,15'd13491,15'd13492,15'd13493,15'd13494,15'd13495,15'd13496,15'd13497,15'd13498,15'd13499,15'd13500,15'd13501,15'd13502,15'd13503,15'd13504,15'd13505,15'd13506,15'd13507,15'd13508,15'd13509,15'd13510,15'd13511,15'd13512,15'd13513,15'd13514,15'd13515,15'd13516,15'd13517,15'd13518,15'd13519,
15'd13760,15'd13761,15'd13762,15'd13763,15'd13764,15'd13765,15'd13766,15'd13767,15'd13768,15'd13769,15'd13770,15'd13771,15'd13772,15'd13773,15'd13774,15'd13775,15'd13776,15'd13777,15'd13778,15'd13779,15'd13780,15'd13781,15'd13782,15'd13783,15'd13784,15'd13785,15'd13786,15'd13787,15'd13788,15'd13789,15'd13790,15'd13791,15'd13792,15'd13793,15'd13794,15'd13795,15'd13796,15'd13797,15'd13798,15'd13799,15'd13800,15'd13801,15'd13802,15'd13803,15'd13804,15'd13805,15'd13806,15'd13807,15'd13808,15'd13809,15'd13810,15'd13811,15'd13812,15'd13813,15'd13814,15'd13815,15'd13816,15'd13817,15'd13818,15'd13819,15'd13820,15'd13821,15'd13822,15'd13823,15'd13824,15'd13825,15'd13826,15'd13827,15'd13828,15'd13829,15'd13830,15'd13831,15'd13832,15'd13833,15'd13834,15'd13835,15'd13836,15'd13837,15'd13838,15'd13839,
15'd14080,15'd14081,15'd14082,15'd14083,15'd14084,15'd14085,15'd14086,15'd14087,15'd14088,15'd14089,15'd14090,15'd14091,15'd14092,15'd14093,15'd14094,15'd14095,15'd14096,15'd14097,15'd14098,15'd14099,15'd14100,15'd14101,15'd14102,15'd14103,15'd14104,15'd14105,15'd14106,15'd14107,15'd14108,15'd14109,15'd14110,15'd14111,15'd14112,15'd14113,15'd14114,15'd14115,15'd14116,15'd14117,15'd14118,15'd14119,15'd14120,15'd14121,15'd14122,15'd14123,15'd14124,15'd14125,15'd14126,15'd14127,15'd14128,15'd14129,15'd14130,15'd14131,15'd14132,15'd14133,15'd14134,15'd14135,15'd14136,15'd14137,15'd14138,15'd14139,15'd14140,15'd14141,15'd14142,15'd14143,15'd14144,15'd14145,15'd14146,15'd14147,15'd14148,15'd14149,15'd14150,15'd14151,15'd14152,15'd14153,15'd14154,15'd14155,15'd14156,15'd14157,15'd14158,15'd14159,
15'd14400,15'd14401,15'd14402,15'd14403,15'd14404,15'd14405,15'd14406,15'd14407,15'd14408,15'd14409,15'd14410,15'd14411,15'd14412,15'd14413,15'd14414,15'd14415,15'd14416,15'd14417,15'd14418,15'd14419,15'd14420,15'd14421,15'd14422,15'd14423,15'd14424,15'd14425,15'd14426,15'd14427,15'd14428,15'd14429,15'd14430,15'd14431,15'd14432,15'd14433,15'd14434,15'd14435,15'd14436,15'd14437,15'd14438,15'd14439,15'd14440,15'd14441,15'd14442,15'd14443,15'd14444,15'd14445,15'd14446,15'd14447,15'd14448,15'd14449,15'd14450,15'd14451,15'd14452,15'd14453,15'd14454,15'd14455,15'd14456,15'd14457,15'd14458,15'd14459,15'd14460,15'd14461,15'd14462,15'd14463,15'd14464,15'd14465,15'd14466,15'd14467,15'd14468,15'd14469,15'd14470,15'd14471,15'd14472,15'd14473,15'd14474,15'd14475,15'd14476,15'd14477,15'd14478,15'd14479,
15'd14720,15'd14721,15'd14722,15'd14723,15'd14724,15'd14725,15'd14726,15'd14727,15'd14728,15'd14729,15'd14730,15'd14731,15'd14732,15'd14733,15'd14734,15'd14735,15'd14736,15'd14737,15'd14738,15'd14739,15'd14740,15'd14741,15'd14742,15'd14743,15'd14744,15'd14745,15'd14746,15'd14747,15'd14748,15'd14749,15'd14750,15'd14751,15'd14752,15'd14753,15'd14754,15'd14755,15'd14756,15'd14757,15'd14758,15'd14759,15'd14760,15'd14761,15'd14762,15'd14763,15'd14764,15'd14765,15'd14766,15'd14767,15'd14768,15'd14769,15'd14770,15'd14771,15'd14772,15'd14773,15'd14774,15'd14775,15'd14776,15'd14777,15'd14778,15'd14779,15'd14780,15'd14781,15'd14782,15'd14783,15'd14784,15'd14785,15'd14786,15'd14787,15'd14788,15'd14789,15'd14790,15'd14791,15'd14792,15'd14793,15'd14794,15'd14795,15'd14796,15'd14797,15'd14798,15'd14799,
15'd15040,15'd15041,15'd15042,15'd15043,15'd15044,15'd15045,15'd15046,15'd15047,15'd15048,15'd15049,15'd15050,15'd15051,15'd15052,15'd15053,15'd15054,15'd15055,15'd15056,15'd15057,15'd15058,15'd15059,15'd15060,15'd15061,15'd15062,15'd15063,15'd15064,15'd15065,15'd15066,15'd15067,15'd15068,15'd15069,15'd15070,15'd15071,15'd15072,15'd15073,15'd15074,15'd15075,15'd15076,15'd15077,15'd15078,15'd15079,15'd15080,15'd15081,15'd15082,15'd15083,15'd15084,15'd15085,15'd15086,15'd15087,15'd15088,15'd15089,15'd15090,15'd15091,15'd15092,15'd15093,15'd15094,15'd15095,15'd15096,15'd15097,15'd15098,15'd15099,15'd15100,15'd15101,15'd15102,15'd15103,15'd15104,15'd15105,15'd15106,15'd15107,15'd15108,15'd15109,15'd15110,15'd15111,15'd15112,15'd15113,15'd15114,15'd15115,15'd15116,15'd15117,15'd15118,15'd15119,
15'd15360,15'd15361,15'd15362,15'd15363,15'd15364,15'd15365,15'd15366,15'd15367,15'd15368,15'd15369,15'd15370,15'd15371,15'd15372,15'd15373,15'd15374,15'd15375,15'd15376,15'd15377,15'd15378,15'd15379,15'd15380,15'd15381,15'd15382,15'd15383,15'd15384,15'd15385,15'd15386,15'd15387,15'd15388,15'd15389,15'd15390,15'd15391,15'd15392,15'd15393,15'd15394,15'd15395,15'd15396,15'd15397,15'd15398,15'd15399,15'd15400,15'd15401,15'd15402,15'd15403,15'd15404,15'd15405,15'd15406,15'd15407,15'd15408,15'd15409,15'd15410,15'd15411,15'd15412,15'd15413,15'd15414,15'd15415,15'd15416,15'd15417,15'd15418,15'd15419,15'd15420,15'd15421,15'd15422,15'd15423,15'd15424,15'd15425,15'd15426,15'd15427,15'd15428,15'd15429,15'd15430,15'd15431,15'd15432,15'd15433,15'd15434,15'd15435,15'd15436,15'd15437,15'd15438,15'd15439,
15'd15680,15'd15681,15'd15682,15'd15683,15'd15684,15'd15685,15'd15686,15'd15687,15'd15688,15'd15689,15'd15690,15'd15691,15'd15692,15'd15693,15'd15694,15'd15695,15'd15696,15'd15697,15'd15698,15'd15699,15'd15700,15'd15701,15'd15702,15'd15703,15'd15704,15'd15705,15'd15706,15'd15707,15'd15708,15'd15709,15'd15710,15'd15711,15'd15712,15'd15713,15'd15714,15'd15715,15'd15716,15'd15717,15'd15718,15'd15719,15'd15720,15'd15721,15'd15722,15'd15723,15'd15724,15'd15725,15'd15726,15'd15727,15'd15728,15'd15729,15'd15730,15'd15731,15'd15732,15'd15733,15'd15734,15'd15735,15'd15736,15'd15737,15'd15738,15'd15739,15'd15740,15'd15741,15'd15742,15'd15743,15'd15744,15'd15745,15'd15746,15'd15747,15'd15748,15'd15749,15'd15750,15'd15751,15'd15752,15'd15753,15'd15754,15'd15755,15'd15756,15'd15757,15'd15758,15'd15759,
15'd16000,15'd16001,15'd16002,15'd16003,15'd16004,15'd16005,15'd16006,15'd16007,15'd16008,15'd16009,15'd16010,15'd16011,15'd16012,15'd16013,15'd16014,15'd16015,15'd16016,15'd16017,15'd16018,15'd16019,15'd16020,15'd16021,15'd16022,15'd16023,15'd16024,15'd16025,15'd16026,15'd16027,15'd16028,15'd16029,15'd16030,15'd16031,15'd16032,15'd16033,15'd16034,15'd16035,15'd16036,15'd16037,15'd16038,15'd16039,15'd16040,15'd16041,15'd16042,15'd16043,15'd16044,15'd16045,15'd16046,15'd16047,15'd16048,15'd16049,15'd16050,15'd16051,15'd16052,15'd16053,15'd16054,15'd16055,15'd16056,15'd16057,15'd16058,15'd16059,15'd16060,15'd16061,15'd16062,15'd16063,15'd16064,15'd16065,15'd16066,15'd16067,15'd16068,15'd16069,15'd16070,15'd16071,15'd16072,15'd16073,15'd16074,15'd16075,15'd16076,15'd16077,15'd16078,15'd16079,
15'd16320,15'd16321,15'd16322,15'd16323,15'd16324,15'd16325,15'd16326,15'd16327,15'd16328,15'd16329,15'd16330,15'd16331,15'd16332,15'd16333,15'd16334,15'd16335,15'd16336,15'd16337,15'd16338,15'd16339,15'd16340,15'd16341,15'd16342,15'd16343,15'd16344,15'd16345,15'd16346,15'd16347,15'd16348,15'd16349,15'd16350,15'd16351,15'd16352,15'd16353,15'd16354,15'd16355,15'd16356,15'd16357,15'd16358,15'd16359,15'd16360,15'd16361,15'd16362,15'd16363,15'd16364,15'd16365,15'd16366,15'd16367,15'd16368,15'd16369,15'd16370,15'd16371,15'd16372,15'd16373,15'd16374,15'd16375,15'd16376,15'd16377,15'd16378,15'd16379,15'd16380,15'd16381,15'd16382,15'd16383,15'd16384,15'd16385,15'd16386,15'd16387,15'd16388,15'd16389,15'd16390,15'd16391,15'd16392,15'd16393,15'd16394,15'd16395,15'd16396,15'd16397,15'd16398,15'd16399,
15'd16640,15'd16641,15'd16642,15'd16643,15'd16644,15'd16645,15'd16646,15'd16647,15'd16648,15'd16649,15'd16650,15'd16651,15'd16652,15'd16653,15'd16654,15'd16655,15'd16656,15'd16657,15'd16658,15'd16659,15'd16660,15'd16661,15'd16662,15'd16663,15'd16664,15'd16665,15'd16666,15'd16667,15'd16668,15'd16669,15'd16670,15'd16671,15'd16672,15'd16673,15'd16674,15'd16675,15'd16676,15'd16677,15'd16678,15'd16679,15'd16680,15'd16681,15'd16682,15'd16683,15'd16684,15'd16685,15'd16686,15'd16687,15'd16688,15'd16689,15'd16690,15'd16691,15'd16692,15'd16693,15'd16694,15'd16695,15'd16696,15'd16697,15'd16698,15'd16699,15'd16700,15'd16701,15'd16702,15'd16703,15'd16704,15'd16705,15'd16706,15'd16707,15'd16708,15'd16709,15'd16710,15'd16711,15'd16712,15'd16713,15'd16714,15'd16715,15'd16716,15'd16717,15'd16718,15'd16719,
15'd16960,15'd16961,15'd16962,15'd16963,15'd16964,15'd16965,15'd16966,15'd16967,15'd16968,15'd16969,15'd16970,15'd16971,15'd16972,15'd16973,15'd16974,15'd16975,15'd16976,15'd16977,15'd16978,15'd16979,15'd16980,15'd16981,15'd16982,15'd16983,15'd16984,15'd16985,15'd16986,15'd16987,15'd16988,15'd16989,15'd16990,15'd16991,15'd16992,15'd16993,15'd16994,15'd16995,15'd16996,15'd16997,15'd16998,15'd16999,15'd17000,15'd17001,15'd17002,15'd17003,15'd17004,15'd17005,15'd17006,15'd17007,15'd17008,15'd17009,15'd17010,15'd17011,15'd17012,15'd17013,15'd17014,15'd17015,15'd17016,15'd17017,15'd17018,15'd17019,15'd17020,15'd17021,15'd17022,15'd17023,15'd17024,15'd17025,15'd17026,15'd17027,15'd17028,15'd17029,15'd17030,15'd17031,15'd17032,15'd17033,15'd17034,15'd17035,15'd17036,15'd17037,15'd17038,15'd17039,
15'd17280,15'd17281,15'd17282,15'd17283,15'd17284,15'd17285,15'd17286,15'd17287,15'd17288,15'd17289,15'd17290,15'd17291,15'd17292,15'd17293,15'd17294,15'd17295,15'd17296,15'd17297,15'd17298,15'd17299,15'd17300,15'd17301,15'd17302,15'd17303,15'd17304,15'd17305,15'd17306,15'd17307,15'd17308,15'd17309,15'd17310,15'd17311,15'd17312,15'd17313,15'd17314,15'd17315,15'd17316,15'd17317,15'd17318,15'd17319,15'd17320,15'd17321,15'd17322,15'd17323,15'd17324,15'd17325,15'd17326,15'd17327,15'd17328,15'd17329,15'd17330,15'd17331,15'd17332,15'd17333,15'd17334,15'd17335,15'd17336,15'd17337,15'd17338,15'd17339,15'd17340,15'd17341,15'd17342,15'd17343,15'd17344,15'd17345,15'd17346,15'd17347,15'd17348,15'd17349,15'd17350,15'd17351,15'd17352,15'd17353,15'd17354,15'd17355,15'd17356,15'd17357,15'd17358,15'd17359,
15'd17600,15'd17601,15'd17602,15'd17603,15'd17604,15'd17605,15'd17606,15'd17607,15'd17608,15'd17609,15'd17610,15'd17611,15'd17612,15'd17613,15'd17614,15'd17615,15'd17616,15'd17617,15'd17618,15'd17619,15'd17620,15'd17621,15'd17622,15'd17623,15'd17624,15'd17625,15'd17626,15'd17627,15'd17628,15'd17629,15'd17630,15'd17631,15'd17632,15'd17633,15'd17634,15'd17635,15'd17636,15'd17637,15'd17638,15'd17639,15'd17640,15'd17641,15'd17642,15'd17643,15'd17644,15'd17645,15'd17646,15'd17647,15'd17648,15'd17649,15'd17650,15'd17651,15'd17652,15'd17653,15'd17654,15'd17655,15'd17656,15'd17657,15'd17658,15'd17659,15'd17660,15'd17661,15'd17662,15'd17663,15'd17664,15'd17665,15'd17666,15'd17667,15'd17668,15'd17669,15'd17670,15'd17671,15'd17672,15'd17673,15'd17674,15'd17675,15'd17676,15'd17677,15'd17678,15'd17679,
15'd17920,15'd17921,15'd17922,15'd17923,15'd17924,15'd17925,15'd17926,15'd17927,15'd17928,15'd17929,15'd17930,15'd17931,15'd17932,15'd17933,15'd17934,15'd17935,15'd17936,15'd17937,15'd17938,15'd17939,15'd17940,15'd17941,15'd17942,15'd17943,15'd17944,15'd17945,15'd17946,15'd17947,15'd17948,15'd17949,15'd17950,15'd17951,15'd17952,15'd17953,15'd17954,15'd17955,15'd17956,15'd17957,15'd17958,15'd17959,15'd17960,15'd17961,15'd17962,15'd17963,15'd17964,15'd17965,15'd17966,15'd17967,15'd17968,15'd17969,15'd17970,15'd17971,15'd17972,15'd17973,15'd17974,15'd17975,15'd17976,15'd17977,15'd17978,15'd17979,15'd17980,15'd17981,15'd17982,15'd17983,15'd17984,15'd17985,15'd17986,15'd17987,15'd17988,15'd17989,15'd17990,15'd17991,15'd17992,15'd17993,15'd17994,15'd17995,15'd17996,15'd17997,15'd17998,15'd17999,
15'd18240,15'd18241,15'd18242,15'd18243,15'd18244,15'd18245,15'd18246,15'd18247,15'd18248,15'd18249,15'd18250,15'd18251,15'd18252,15'd18253,15'd18254,15'd18255,15'd18256,15'd18257,15'd18258,15'd18259,15'd18260,15'd18261,15'd18262,15'd18263,15'd18264,15'd18265,15'd18266,15'd18267,15'd18268,15'd18269,15'd18270,15'd18271,15'd18272,15'd18273,15'd18274,15'd18275,15'd18276,15'd18277,15'd18278,15'd18279,15'd18280,15'd18281,15'd18282,15'd18283,15'd18284,15'd18285,15'd18286,15'd18287,15'd18288,15'd18289,15'd18290,15'd18291,15'd18292,15'd18293,15'd18294,15'd18295,15'd18296,15'd18297,15'd18298,15'd18299,15'd18300,15'd18301,15'd18302,15'd18303,15'd18304,15'd18305,15'd18306,15'd18307,15'd18308,15'd18309,15'd18310,15'd18311,15'd18312,15'd18313,15'd18314,15'd18315,15'd18316,15'd18317,15'd18318,15'd18319,
15'd18560,15'd18561,15'd18562,15'd18563,15'd18564,15'd18565,15'd18566,15'd18567,15'd18568,15'd18569,15'd18570,15'd18571,15'd18572,15'd18573,15'd18574,15'd18575,15'd18576,15'd18577,15'd18578,15'd18579,15'd18580,15'd18581,15'd18582,15'd18583,15'd18584,15'd18585,15'd18586,15'd18587,15'd18588,15'd18589,15'd18590,15'd18591,15'd18592,15'd18593,15'd18594,15'd18595,15'd18596,15'd18597,15'd18598,15'd18599,15'd18600,15'd18601,15'd18602,15'd18603,15'd18604,15'd18605,15'd18606,15'd18607,15'd18608,15'd18609,15'd18610,15'd18611,15'd18612,15'd18613,15'd18614,15'd18615,15'd18616,15'd18617,15'd18618,15'd18619,15'd18620,15'd18621,15'd18622,15'd18623,15'd18624,15'd18625,15'd18626,15'd18627,15'd18628,15'd18629,15'd18630,15'd18631,15'd18632,15'd18633,15'd18634,15'd18635,15'd18636,15'd18637,15'd18638,15'd18639,
15'd18880,15'd18881,15'd18882,15'd18883,15'd18884,15'd18885,15'd18886,15'd18887,15'd18888,15'd18889,15'd18890,15'd18891,15'd18892,15'd18893,15'd18894,15'd18895,15'd18896,15'd18897,15'd18898,15'd18899,15'd18900,15'd18901,15'd18902,15'd18903,15'd18904,15'd18905,15'd18906,15'd18907,15'd18908,15'd18909,15'd18910,15'd18911,15'd18912,15'd18913,15'd18914,15'd18915,15'd18916,15'd18917,15'd18918,15'd18919,15'd18920,15'd18921,15'd18922,15'd18923,15'd18924,15'd18925,15'd18926,15'd18927,15'd18928,15'd18929,15'd18930,15'd18931,15'd18932,15'd18933,15'd18934,15'd18935,15'd18936,15'd18937,15'd18938,15'd18939,15'd18940,15'd18941,15'd18942,15'd18943,15'd18944,15'd18945,15'd18946,15'd18947,15'd18948,15'd18949,15'd18950,15'd18951,15'd18952,15'd18953,15'd18954,15'd18955,15'd18956,15'd18957,15'd18958,15'd18959,
15'd19200,15'd19201,15'd19202,15'd19203,15'd19204,15'd19205,15'd19206,15'd19207,15'd19208,15'd19209,15'd19210,15'd19211,15'd19212,15'd19213,15'd19214,15'd19215,15'd19216,15'd19217,15'd19218,15'd19219,15'd19220,15'd19221,15'd19222,15'd19223,15'd19224,15'd19225,15'd19226,15'd19227,15'd19228,15'd19229,15'd19230,15'd19231,15'd19232,15'd19233,15'd19234,15'd19235,15'd19236,15'd19237,15'd19238,15'd19239,15'd19240,15'd19241,15'd19242,15'd19243,15'd19244,15'd19245,15'd19246,15'd19247,15'd19248,15'd19249,15'd19250,15'd19251,15'd19252,15'd19253,15'd19254,15'd19255,15'd19256,15'd19257,15'd19258,15'd19259,15'd19260,15'd19261,15'd19262,15'd19263,15'd19264,15'd19265,15'd19266,15'd19267,15'd19268,15'd19269,15'd19270,15'd19271,15'd19272,15'd19273,15'd19274,15'd19275,15'd19276,15'd19277,15'd19278,15'd19279,
15'd19520,15'd19521,15'd19522,15'd19523,15'd19524,15'd19525,15'd19526,15'd19527,15'd19528,15'd19529,15'd19530,15'd19531,15'd19532,15'd19533,15'd19534,15'd19535,15'd19536,15'd19537,15'd19538,15'd19539,15'd19540,15'd19541,15'd19542,15'd19543,15'd19544,15'd19545,15'd19546,15'd19547,15'd19548,15'd19549,15'd19550,15'd19551,15'd19552,15'd19553,15'd19554,15'd19555,15'd19556,15'd19557,15'd19558,15'd19559,15'd19560,15'd19561,15'd19562,15'd19563,15'd19564,15'd19565,15'd19566,15'd19567,15'd19568,15'd19569,15'd19570,15'd19571,15'd19572,15'd19573,15'd19574,15'd19575,15'd19576,15'd19577,15'd19578,15'd19579,15'd19580,15'd19581,15'd19582,15'd19583,15'd19584,15'd19585,15'd19586,15'd19587,15'd19588,15'd19589,15'd19590,15'd19591,15'd19592,15'd19593,15'd19594,15'd19595,15'd19596,15'd19597,15'd19598,15'd19599,
15'd19840,15'd19841,15'd19842,15'd19843,15'd19844,15'd19845,15'd19846,15'd19847,15'd19848,15'd19849,15'd19850,15'd19851,15'd19852,15'd19853,15'd19854,15'd19855,15'd19856,15'd19857,15'd19858,15'd19859,15'd19860,15'd19861,15'd19862,15'd19863,15'd19864,15'd19865,15'd19866,15'd19867,15'd19868,15'd19869,15'd19870,15'd19871,15'd19872,15'd19873,15'd19874,15'd19875,15'd19876,15'd19877,15'd19878,15'd19879,15'd19880,15'd19881,15'd19882,15'd19883,15'd19884,15'd19885,15'd19886,15'd19887,15'd19888,15'd19889,15'd19890,15'd19891,15'd19892,15'd19893,15'd19894,15'd19895,15'd19896,15'd19897,15'd19898,15'd19899,15'd19900,15'd19901,15'd19902,15'd19903,15'd19904,15'd19905,15'd19906,15'd19907,15'd19908,15'd19909,15'd19910,15'd19911,15'd19912,15'd19913,15'd19914,15'd19915,15'd19916,15'd19917,15'd19918,15'd19919,
15'd20160,15'd20161,15'd20162,15'd20163,15'd20164,15'd20165,15'd20166,15'd20167,15'd20168,15'd20169,15'd20170,15'd20171,15'd20172,15'd20173,15'd20174,15'd20175,15'd20176,15'd20177,15'd20178,15'd20179,15'd20180,15'd20181,15'd20182,15'd20183,15'd20184,15'd20185,15'd20186,15'd20187,15'd20188,15'd20189,15'd20190,15'd20191,15'd20192,15'd20193,15'd20194,15'd20195,15'd20196,15'd20197,15'd20198,15'd20199,15'd20200,15'd20201,15'd20202,15'd20203,15'd20204,15'd20205,15'd20206,15'd20207,15'd20208,15'd20209,15'd20210,15'd20211,15'd20212,15'd20213,15'd20214,15'd20215,15'd20216,15'd20217,15'd20218,15'd20219,15'd20220,15'd20221,15'd20222,15'd20223,15'd20224,15'd20225,15'd20226,15'd20227,15'd20228,15'd20229,15'd20230,15'd20231,15'd20232,15'd20233,15'd20234,15'd20235,15'd20236,15'd20237,15'd20238,15'd20239,
15'd20480,15'd20481,15'd20482,15'd20483,15'd20484,15'd20485,15'd20486,15'd20487,15'd20488,15'd20489,15'd20490,15'd20491,15'd20492,15'd20493,15'd20494,15'd20495,15'd20496,15'd20497,15'd20498,15'd20499,15'd20500,15'd20501,15'd20502,15'd20503,15'd20504,15'd20505,15'd20506,15'd20507,15'd20508,15'd20509,15'd20510,15'd20511,15'd20512,15'd20513,15'd20514,15'd20515,15'd20516,15'd20517,15'd20518,15'd20519,15'd20520,15'd20521,15'd20522,15'd20523,15'd20524,15'd20525,15'd20526,15'd20527,15'd20528,15'd20529,15'd20530,15'd20531,15'd20532,15'd20533,15'd20534,15'd20535,15'd20536,15'd20537,15'd20538,15'd20539,15'd20540,15'd20541,15'd20542,15'd20543,15'd20544,15'd20545,15'd20546,15'd20547,15'd20548,15'd20549,15'd20550,15'd20551,15'd20552,15'd20553,15'd20554,15'd20555,15'd20556,15'd20557,15'd20558,15'd20559,
15'd20800,15'd20801,15'd20802,15'd20803,15'd20804,15'd20805,15'd20806,15'd20807,15'd20808,15'd20809,15'd20810,15'd20811,15'd20812,15'd20813,15'd20814,15'd20815,15'd20816,15'd20817,15'd20818,15'd20819,15'd20820,15'd20821,15'd20822,15'd20823,15'd20824,15'd20825,15'd20826,15'd20827,15'd20828,15'd20829,15'd20830,15'd20831,15'd20832,15'd20833,15'd20834,15'd20835,15'd20836,15'd20837,15'd20838,15'd20839,15'd20840,15'd20841,15'd20842,15'd20843,15'd20844,15'd20845,15'd20846,15'd20847,15'd20848,15'd20849,15'd20850,15'd20851,15'd20852,15'd20853,15'd20854,15'd20855,15'd20856,15'd20857,15'd20858,15'd20859,15'd20860,15'd20861,15'd20862,15'd20863,15'd20864,15'd20865,15'd20866,15'd20867,15'd20868,15'd20869,15'd20870,15'd20871,15'd20872,15'd20873,15'd20874,15'd20875,15'd20876,15'd20877,15'd20878,15'd20879,
15'd21120,15'd21121,15'd21122,15'd21123,15'd21124,15'd21125,15'd21126,15'd21127,15'd21128,15'd21129,15'd21130,15'd21131,15'd21132,15'd21133,15'd21134,15'd21135,15'd21136,15'd21137,15'd21138,15'd21139,15'd21140,15'd21141,15'd21142,15'd21143,15'd21144,15'd21145,15'd21146,15'd21147,15'd21148,15'd21149,15'd21150,15'd21151,15'd21152,15'd21153,15'd21154,15'd21155,15'd21156,15'd21157,15'd21158,15'd21159,15'd21160,15'd21161,15'd21162,15'd21163,15'd21164,15'd21165,15'd21166,15'd21167,15'd21168,15'd21169,15'd21170,15'd21171,15'd21172,15'd21173,15'd21174,15'd21175,15'd21176,15'd21177,15'd21178,15'd21179,15'd21180,15'd21181,15'd21182,15'd21183,15'd21184,15'd21185,15'd21186,15'd21187,15'd21188,15'd21189,15'd21190,15'd21191,15'd21192,15'd21193,15'd21194,15'd21195,15'd21196,15'd21197,15'd21198,15'd21199,
15'd21440,15'd21441,15'd21442,15'd21443,15'd21444,15'd21445,15'd21446,15'd21447,15'd21448,15'd21449,15'd21450,15'd21451,15'd21452,15'd21453,15'd21454,15'd21455,15'd21456,15'd21457,15'd21458,15'd21459,15'd21460,15'd21461,15'd21462,15'd21463,15'd21464,15'd21465,15'd21466,15'd21467,15'd21468,15'd21469,15'd21470,15'd21471,15'd21472,15'd21473,15'd21474,15'd21475,15'd21476,15'd21477,15'd21478,15'd21479,15'd21480,15'd21481,15'd21482,15'd21483,15'd21484,15'd21485,15'd21486,15'd21487,15'd21488,15'd21489,15'd21490,15'd21491,15'd21492,15'd21493,15'd21494,15'd21495,15'd21496,15'd21497,15'd21498,15'd21499,15'd21500,15'd21501,15'd21502,15'd21503,15'd21504,15'd21505,15'd21506,15'd21507,15'd21508,15'd21509,15'd21510,15'd21511,15'd21512,15'd21513,15'd21514,15'd21515,15'd21516,15'd21517,15'd21518,15'd21519,
15'd21760,15'd21761,15'd21762,15'd21763,15'd21764,15'd21765,15'd21766,15'd21767,15'd21768,15'd21769,15'd21770,15'd21771,15'd21772,15'd21773,15'd21774,15'd21775,15'd21776,15'd21777,15'd21778,15'd21779,15'd21780,15'd21781,15'd21782,15'd21783,15'd21784,15'd21785,15'd21786,15'd21787,15'd21788,15'd21789,15'd21790,15'd21791,15'd21792,15'd21793,15'd21794,15'd21795,15'd21796,15'd21797,15'd21798,15'd21799,15'd21800,15'd21801,15'd21802,15'd21803,15'd21804,15'd21805,15'd21806,15'd21807,15'd21808,15'd21809,15'd21810,15'd21811,15'd21812,15'd21813,15'd21814,15'd21815,15'd21816,15'd21817,15'd21818,15'd21819,15'd21820,15'd21821,15'd21822,15'd21823,15'd21824,15'd21825,15'd21826,15'd21827,15'd21828,15'd21829,15'd21830,15'd21831,15'd21832,15'd21833,15'd21834,15'd21835,15'd21836,15'd21837,15'd21838,15'd21839,
15'd22080,15'd22081,15'd22082,15'd22083,15'd22084,15'd22085,15'd22086,15'd22087,15'd22088,15'd22089,15'd22090,15'd22091,15'd22092,15'd22093,15'd22094,15'd22095,15'd22096,15'd22097,15'd22098,15'd22099,15'd22100,15'd22101,15'd22102,15'd22103,15'd22104,15'd22105,15'd22106,15'd22107,15'd22108,15'd22109,15'd22110,15'd22111,15'd22112,15'd22113,15'd22114,15'd22115,15'd22116,15'd22117,15'd22118,15'd22119,15'd22120,15'd22121,15'd22122,15'd22123,15'd22124,15'd22125,15'd22126,15'd22127,15'd22128,15'd22129,15'd22130,15'd22131,15'd22132,15'd22133,15'd22134,15'd22135,15'd22136,15'd22137,15'd22138,15'd22139,15'd22140,15'd22141,15'd22142,15'd22143,15'd22144,15'd22145,15'd22146,15'd22147,15'd22148,15'd22149,15'd22150,15'd22151,15'd22152,15'd22153,15'd22154,15'd22155,15'd22156,15'd22157,15'd22158,15'd22159,
15'd22400,15'd22401,15'd22402,15'd22403,15'd22404,15'd22405,15'd22406,15'd22407,15'd22408,15'd22409,15'd22410,15'd22411,15'd22412,15'd22413,15'd22414,15'd22415,15'd22416,15'd22417,15'd22418,15'd22419,15'd22420,15'd22421,15'd22422,15'd22423,15'd22424,15'd22425,15'd22426,15'd22427,15'd22428,15'd22429,15'd22430,15'd22431,15'd22432,15'd22433,15'd22434,15'd22435,15'd22436,15'd22437,15'd22438,15'd22439,15'd22440,15'd22441,15'd22442,15'd22443,15'd22444,15'd22445,15'd22446,15'd22447,15'd22448,15'd22449,15'd22450,15'd22451,15'd22452,15'd22453,15'd22454,15'd22455,15'd22456,15'd22457,15'd22458,15'd22459,15'd22460,15'd22461,15'd22462,15'd22463,15'd22464,15'd22465,15'd22466,15'd22467,15'd22468,15'd22469,15'd22470,15'd22471,15'd22472,15'd22473,15'd22474,15'd22475,15'd22476,15'd22477,15'd22478,15'd22479,
15'd22720,15'd22721,15'd22722,15'd22723,15'd22724,15'd22725,15'd22726,15'd22727,15'd22728,15'd22729,15'd22730,15'd22731,15'd22732,15'd22733,15'd22734,15'd22735,15'd22736,15'd22737,15'd22738,15'd22739,15'd22740,15'd22741,15'd22742,15'd22743,15'd22744,15'd22745,15'd22746,15'd22747,15'd22748,15'd22749,15'd22750,15'd22751,15'd22752,15'd22753,15'd22754,15'd22755,15'd22756,15'd22757,15'd22758,15'd22759,15'd22760,15'd22761,15'd22762,15'd22763,15'd22764,15'd22765,15'd22766,15'd22767,15'd22768,15'd22769,15'd22770,15'd22771,15'd22772,15'd22773,15'd22774,15'd22775,15'd22776,15'd22777,15'd22778,15'd22779,15'd22780,15'd22781,15'd22782,15'd22783,15'd22784,15'd22785,15'd22786,15'd22787,15'd22788,15'd22789,15'd22790,15'd22791,15'd22792,15'd22793,15'd22794,15'd22795,15'd22796,15'd22797,15'd22798,15'd22799,
15'd23040,15'd23041,15'd23042,15'd23043,15'd23044,15'd23045,15'd23046,15'd23047,15'd23048,15'd23049,15'd23050,15'd23051,15'd23052,15'd23053,15'd23054,15'd23055,15'd23056,15'd23057,15'd23058,15'd23059,15'd23060,15'd23061,15'd23062,15'd23063,15'd23064,15'd23065,15'd23066,15'd23067,15'd23068,15'd23069,15'd23070,15'd23071,15'd23072,15'd23073,15'd23074,15'd23075,15'd23076,15'd23077,15'd23078,15'd23079,15'd23080,15'd23081,15'd23082,15'd23083,15'd23084,15'd23085,15'd23086,15'd23087,15'd23088,15'd23089,15'd23090,15'd23091,15'd23092,15'd23093,15'd23094,15'd23095,15'd23096,15'd23097,15'd23098,15'd23099,15'd23100,15'd23101,15'd23102,15'd23103,15'd23104,15'd23105,15'd23106,15'd23107,15'd23108,15'd23109,15'd23110,15'd23111,15'd23112,15'd23113,15'd23114,15'd23115,15'd23116,15'd23117,15'd23118,15'd23119,
15'd23360,15'd23361,15'd23362,15'd23363,15'd23364,15'd23365,15'd23366,15'd23367,15'd23368,15'd23369,15'd23370,15'd23371,15'd23372,15'd23373,15'd23374,15'd23375,15'd23376,15'd23377,15'd23378,15'd23379,15'd23380,15'd23381,15'd23382,15'd23383,15'd23384,15'd23385,15'd23386,15'd23387,15'd23388,15'd23389,15'd23390,15'd23391,15'd23392,15'd23393,15'd23394,15'd23395,15'd23396,15'd23397,15'd23398,15'd23399,15'd23400,15'd23401,15'd23402,15'd23403,15'd23404,15'd23405,15'd23406,15'd23407,15'd23408,15'd23409,15'd23410,15'd23411,15'd23412,15'd23413,15'd23414,15'd23415,15'd23416,15'd23417,15'd23418,15'd23419,15'd23420,15'd23421,15'd23422,15'd23423,15'd23424,15'd23425,15'd23426,15'd23427,15'd23428,15'd23429,15'd23430,15'd23431,15'd23432,15'd23433,15'd23434,15'd23435,15'd23436,15'd23437,15'd23438,15'd23439,
15'd23680,15'd23681,15'd23682,15'd23683,15'd23684,15'd23685,15'd23686,15'd23687,15'd23688,15'd23689,15'd23690,15'd23691,15'd23692,15'd23693,15'd23694,15'd23695,15'd23696,15'd23697,15'd23698,15'd23699,15'd23700,15'd23701,15'd23702,15'd23703,15'd23704,15'd23705,15'd23706,15'd23707,15'd23708,15'd23709,15'd23710,15'd23711,15'd23712,15'd23713,15'd23714,15'd23715,15'd23716,15'd23717,15'd23718,15'd23719,15'd23720,15'd23721,15'd23722,15'd23723,15'd23724,15'd23725,15'd23726,15'd23727,15'd23728,15'd23729,15'd23730,15'd23731,15'd23732,15'd23733,15'd23734,15'd23735,15'd23736,15'd23737,15'd23738,15'd23739,15'd23740,15'd23741,15'd23742,15'd23743,15'd23744,15'd23745,15'd23746,15'd23747,15'd23748,15'd23749,15'd23750,15'd23751,15'd23752,15'd23753,15'd23754,15'd23755,15'd23756,15'd23757,15'd23758,15'd23759,
15'd24000,15'd24001,15'd24002,15'd24003,15'd24004,15'd24005,15'd24006,15'd24007,15'd24008,15'd24009,15'd24010,15'd24011,15'd24012,15'd24013,15'd24014,15'd24015,15'd24016,15'd24017,15'd24018,15'd24019,15'd24020,15'd24021,15'd24022,15'd24023,15'd24024,15'd24025,15'd24026,15'd24027,15'd24028,15'd24029,15'd24030,15'd24031,15'd24032,15'd24033,15'd24034,15'd24035,15'd24036,15'd24037,15'd24038,15'd24039,15'd24040,15'd24041,15'd24042,15'd24043,15'd24044,15'd24045,15'd24046,15'd24047,15'd24048,15'd24049,15'd24050,15'd24051,15'd24052,15'd24053,15'd24054,15'd24055,15'd24056,15'd24057,15'd24058,15'd24059,15'd24060,15'd24061,15'd24062,15'd24063,15'd24064,15'd24065,15'd24066,15'd24067,15'd24068,15'd24069,15'd24070,15'd24071,15'd24072,15'd24073,15'd24074,15'd24075,15'd24076,15'd24077,15'd24078,15'd24079,
15'd24320,15'd24321,15'd24322,15'd24323,15'd24324,15'd24325,15'd24326,15'd24327,15'd24328,15'd24329,15'd24330,15'd24331,15'd24332,15'd24333,15'd24334,15'd24335,15'd24336,15'd24337,15'd24338,15'd24339,15'd24340,15'd24341,15'd24342,15'd24343,15'd24344,15'd24345,15'd24346,15'd24347,15'd24348,15'd24349,15'd24350,15'd24351,15'd24352,15'd24353,15'd24354,15'd24355,15'd24356,15'd24357,15'd24358,15'd24359,15'd24360,15'd24361,15'd24362,15'd24363,15'd24364,15'd24365,15'd24366,15'd24367,15'd24368,15'd24369,15'd24370,15'd24371,15'd24372,15'd24373,15'd24374,15'd24375,15'd24376,15'd24377,15'd24378,15'd24379,15'd24380,15'd24381,15'd24382,15'd24383,15'd24384,15'd24385,15'd24386,15'd24387,15'd24388,15'd24389,15'd24390,15'd24391,15'd24392,15'd24393,15'd24394,15'd24395,15'd24396,15'd24397,15'd24398,15'd24399,
15'd24640,15'd24641,15'd24642,15'd24643,15'd24644,15'd24645,15'd24646,15'd24647,15'd24648,15'd24649,15'd24650,15'd24651,15'd24652,15'd24653,15'd24654,15'd24655,15'd24656,15'd24657,15'd24658,15'd24659,15'd24660,15'd24661,15'd24662,15'd24663,15'd24664,15'd24665,15'd24666,15'd24667,15'd24668,15'd24669,15'd24670,15'd24671,15'd24672,15'd24673,15'd24674,15'd24675,15'd24676,15'd24677,15'd24678,15'd24679,15'd24680,15'd24681,15'd24682,15'd24683,15'd24684,15'd24685,15'd24686,15'd24687,15'd24688,15'd24689,15'd24690,15'd24691,15'd24692,15'd24693,15'd24694,15'd24695,15'd24696,15'd24697,15'd24698,15'd24699,15'd24700,15'd24701,15'd24702,15'd24703,15'd24704,15'd24705,15'd24706,15'd24707,15'd24708,15'd24709,15'd24710,15'd24711,15'd24712,15'd24713,15'd24714,15'd24715,15'd24716,15'd24717,15'd24718,15'd24719,
15'd24960,15'd24961,15'd24962,15'd24963,15'd24964,15'd24965,15'd24966,15'd24967,15'd24968,15'd24969,15'd24970,15'd24971,15'd24972,15'd24973,15'd24974,15'd24975,15'd24976,15'd24977,15'd24978,15'd24979,15'd24980,15'd24981,15'd24982,15'd24983,15'd24984,15'd24985,15'd24986,15'd24987,15'd24988,15'd24989,15'd24990,15'd24991,15'd24992,15'd24993,15'd24994,15'd24995,15'd24996,15'd24997,15'd24998,15'd24999,15'd25000,15'd25001,15'd25002,15'd25003,15'd25004,15'd25005,15'd25006,15'd25007,15'd25008,15'd25009,15'd25010,15'd25011,15'd25012,15'd25013,15'd25014,15'd25015,15'd25016,15'd25017,15'd25018,15'd25019,15'd25020,15'd25021,15'd25022,15'd25023,15'd25024,15'd25025,15'd25026,15'd25027,15'd25028,15'd25029,15'd25030,15'd25031,15'd25032,15'd25033,15'd25034,15'd25035,15'd25036,15'd25037,15'd25038,15'd25039,
15'd25280,15'd25281,15'd25282,15'd25283,15'd25284,15'd25285,15'd25286,15'd25287,15'd25288,15'd25289,15'd25290,15'd25291,15'd25292,15'd25293,15'd25294,15'd25295,15'd25296,15'd25297,15'd25298,15'd25299,15'd25300,15'd25301,15'd25302,15'd25303,15'd25304,15'd25305,15'd25306,15'd25307,15'd25308,15'd25309,15'd25310,15'd25311,15'd25312,15'd25313,15'd25314,15'd25315,15'd25316,15'd25317,15'd25318,15'd25319,15'd25320,15'd25321,15'd25322,15'd25323,15'd25324,15'd25325,15'd25326,15'd25327,15'd25328,15'd25329,15'd25330,15'd25331,15'd25332,15'd25333,15'd25334,15'd25335,15'd25336,15'd25337,15'd25338,15'd25339,15'd25340,15'd25341,15'd25342,15'd25343,15'd25344,15'd25345,15'd25346,15'd25347,15'd25348,15'd25349,15'd25350,15'd25351,15'd25352,15'd25353,15'd25354,15'd25355,15'd25356,15'd25357,15'd25358,15'd25359};
parameter [14:0] state_1 [0:6399] = {
15'd25280,15'd24960,15'd24640,15'd24320,15'd24000,15'd23680,15'd23360,15'd23040,15'd22720,15'd22400,15'd22080,15'd21760,15'd21440,15'd21120,15'd20800,15'd20480,15'd20160,15'd19840,15'd19520,15'd19200,15'd18880,15'd18560,15'd18240,15'd17920,15'd17600,15'd17280,15'd16960,15'd16640,15'd16320,15'd16000,15'd15680,15'd15360,15'd15040,15'd14720,15'd14400,15'd14080,15'd13760,15'd13440,15'd13120,15'd12800,15'd12480,15'd12160,15'd11840,15'd11520,15'd11200,15'd10880,15'd10560,15'd10240,15'd9920,15'd9600,15'd9280,15'd8960,15'd8640,15'd8320,15'd8000,15'd7680,15'd7360,15'd7040,15'd6720,15'd6400,15'd6080,15'd5760,15'd5440,15'd5120,15'd4800,15'd4480,15'd4160,15'd3840,15'd3520,15'd3200,15'd2880,15'd2560,15'd2240,15'd1920,15'd1600,15'd1280,15'd960,15'd640,15'd320,15'd0,
15'd25281,15'd24961,15'd24641,15'd24321,15'd24001,15'd23681,15'd23361,15'd23041,15'd22721,15'd22401,15'd22081,15'd21761,15'd21441,15'd21121,15'd20801,15'd20481,15'd20161,15'd19841,15'd19521,15'd19201,15'd18881,15'd18561,15'd18241,15'd17921,15'd17601,15'd17281,15'd16961,15'd16641,15'd16321,15'd16001,15'd15681,15'd15361,15'd15041,15'd14721,15'd14401,15'd14081,15'd13761,15'd13441,15'd13121,15'd12801,15'd12481,15'd12161,15'd11841,15'd11521,15'd11201,15'd10881,15'd10561,15'd10241,15'd9921,15'd9601,15'd9281,15'd8961,15'd8641,15'd8321,15'd8001,15'd7681,15'd7361,15'd7041,15'd6721,15'd6401,15'd6081,15'd5761,15'd5441,15'd5121,15'd4801,15'd4481,15'd4161,15'd3841,15'd3521,15'd3201,15'd2881,15'd2561,15'd2241,15'd1921,15'd1601,15'd1281,15'd961,15'd641,15'd321,15'd1,
15'd25282,15'd24962,15'd24642,15'd24322,15'd24002,15'd23682,15'd23362,15'd23042,15'd22722,15'd22402,15'd22082,15'd21762,15'd21442,15'd21122,15'd20802,15'd20482,15'd20162,15'd19842,15'd19522,15'd19202,15'd18882,15'd18562,15'd18242,15'd17922,15'd17602,15'd17282,15'd16962,15'd16642,15'd16322,15'd16002,15'd15682,15'd15362,15'd15042,15'd14722,15'd14402,15'd14082,15'd13762,15'd13442,15'd13122,15'd12802,15'd12482,15'd12162,15'd11842,15'd11522,15'd11202,15'd10882,15'd10562,15'd10242,15'd9922,15'd9602,15'd9282,15'd8962,15'd8642,15'd8322,15'd8002,15'd7682,15'd7362,15'd7042,15'd6722,15'd6402,15'd6082,15'd5762,15'd5442,15'd5122,15'd4802,15'd4482,15'd4162,15'd3842,15'd3522,15'd3202,15'd2882,15'd2562,15'd2242,15'd1922,15'd1602,15'd1282,15'd962,15'd642,15'd322,15'd2,
15'd25283,15'd24963,15'd24643,15'd24323,15'd24003,15'd23683,15'd23363,15'd23043,15'd22723,15'd22403,15'd22083,15'd21763,15'd21443,15'd21123,15'd20803,15'd20483,15'd20163,15'd19843,15'd19523,15'd19203,15'd18883,15'd18563,15'd18243,15'd17923,15'd17603,15'd17283,15'd16963,15'd16643,15'd16323,15'd16003,15'd15683,15'd15363,15'd15043,15'd14723,15'd14403,15'd14083,15'd13763,15'd13443,15'd13123,15'd12803,15'd12483,15'd12163,15'd11843,15'd11523,15'd11203,15'd10883,15'd10563,15'd10243,15'd9923,15'd9603,15'd9283,15'd8963,15'd8643,15'd8323,15'd8003,15'd7683,15'd7363,15'd7043,15'd6723,15'd6403,15'd6083,15'd5763,15'd5443,15'd5123,15'd4803,15'd4483,15'd4163,15'd3843,15'd3523,15'd3203,15'd2883,15'd2563,15'd2243,15'd1923,15'd1603,15'd1283,15'd963,15'd643,15'd323,15'd3,
15'd25284,15'd24964,15'd24644,15'd24324,15'd24004,15'd23684,15'd23364,15'd23044,15'd22724,15'd22404,15'd22084,15'd21764,15'd21444,15'd21124,15'd20804,15'd20484,15'd20164,15'd19844,15'd19524,15'd19204,15'd18884,15'd18564,15'd18244,15'd17924,15'd17604,15'd17284,15'd16964,15'd16644,15'd16324,15'd16004,15'd15684,15'd15364,15'd15044,15'd14724,15'd14404,15'd14084,15'd13764,15'd13444,15'd13124,15'd12804,15'd12484,15'd12164,15'd11844,15'd11524,15'd11204,15'd10884,15'd10564,15'd10244,15'd9924,15'd9604,15'd9284,15'd8964,15'd8644,15'd8324,15'd8004,15'd7684,15'd7364,15'd7044,15'd6724,15'd6404,15'd6084,15'd5764,15'd5444,15'd5124,15'd4804,15'd4484,15'd4164,15'd3844,15'd3524,15'd3204,15'd2884,15'd2564,15'd2244,15'd1924,15'd1604,15'd1284,15'd964,15'd644,15'd324,15'd4,
15'd25285,15'd24965,15'd24645,15'd24325,15'd24005,15'd23685,15'd23365,15'd23045,15'd22725,15'd22405,15'd22085,15'd21765,15'd21445,15'd21125,15'd20805,15'd20485,15'd20165,15'd19845,15'd19525,15'd19205,15'd18885,15'd18565,15'd18245,15'd17925,15'd17605,15'd17285,15'd16965,15'd16645,15'd16325,15'd16005,15'd15685,15'd15365,15'd15045,15'd14725,15'd14405,15'd14085,15'd13765,15'd13445,15'd13125,15'd12805,15'd12485,15'd12165,15'd11845,15'd11525,15'd11205,15'd10885,15'd10565,15'd10245,15'd9925,15'd9605,15'd9285,15'd8965,15'd8645,15'd8325,15'd8005,15'd7685,15'd7365,15'd7045,15'd6725,15'd6405,15'd6085,15'd5765,15'd5445,15'd5125,15'd4805,15'd4485,15'd4165,15'd3845,15'd3525,15'd3205,15'd2885,15'd2565,15'd2245,15'd1925,15'd1605,15'd1285,15'd965,15'd645,15'd325,15'd5,
15'd25286,15'd24966,15'd24646,15'd24326,15'd24006,15'd23686,15'd23366,15'd23046,15'd22726,15'd22406,15'd22086,15'd21766,15'd21446,15'd21126,15'd20806,15'd20486,15'd20166,15'd19846,15'd19526,15'd19206,15'd18886,15'd18566,15'd18246,15'd17926,15'd17606,15'd17286,15'd16966,15'd16646,15'd16326,15'd16006,15'd15686,15'd15366,15'd15046,15'd14726,15'd14406,15'd14086,15'd13766,15'd13446,15'd13126,15'd12806,15'd12486,15'd12166,15'd11846,15'd11526,15'd11206,15'd10886,15'd10566,15'd10246,15'd9926,15'd9606,15'd9286,15'd8966,15'd8646,15'd8326,15'd8006,15'd7686,15'd7366,15'd7046,15'd6726,15'd6406,15'd6086,15'd5766,15'd5446,15'd5126,15'd4806,15'd4486,15'd4166,15'd3846,15'd3526,15'd3206,15'd2886,15'd2566,15'd2246,15'd1926,15'd1606,15'd1286,15'd966,15'd646,15'd326,15'd6,
15'd25287,15'd24967,15'd24647,15'd24327,15'd24007,15'd23687,15'd23367,15'd23047,15'd22727,15'd22407,15'd22087,15'd21767,15'd21447,15'd21127,15'd20807,15'd20487,15'd20167,15'd19847,15'd19527,15'd19207,15'd18887,15'd18567,15'd18247,15'd17927,15'd17607,15'd17287,15'd16967,15'd16647,15'd16327,15'd16007,15'd15687,15'd15367,15'd15047,15'd14727,15'd14407,15'd14087,15'd13767,15'd13447,15'd13127,15'd12807,15'd12487,15'd12167,15'd11847,15'd11527,15'd11207,15'd10887,15'd10567,15'd10247,15'd9927,15'd9607,15'd9287,15'd8967,15'd8647,15'd8327,15'd8007,15'd7687,15'd7367,15'd7047,15'd6727,15'd6407,15'd6087,15'd5767,15'd5447,15'd5127,15'd4807,15'd4487,15'd4167,15'd3847,15'd3527,15'd3207,15'd2887,15'd2567,15'd2247,15'd1927,15'd1607,15'd1287,15'd967,15'd647,15'd327,15'd7,
15'd25288,15'd24968,15'd24648,15'd24328,15'd24008,15'd23688,15'd23368,15'd23048,15'd22728,15'd22408,15'd22088,15'd21768,15'd21448,15'd21128,15'd20808,15'd20488,15'd20168,15'd19848,15'd19528,15'd19208,15'd18888,15'd18568,15'd18248,15'd17928,15'd17608,15'd17288,15'd16968,15'd16648,15'd16328,15'd16008,15'd15688,15'd15368,15'd15048,15'd14728,15'd14408,15'd14088,15'd13768,15'd13448,15'd13128,15'd12808,15'd12488,15'd12168,15'd11848,15'd11528,15'd11208,15'd10888,15'd10568,15'd10248,15'd9928,15'd9608,15'd9288,15'd8968,15'd8648,15'd8328,15'd8008,15'd7688,15'd7368,15'd7048,15'd6728,15'd6408,15'd6088,15'd5768,15'd5448,15'd5128,15'd4808,15'd4488,15'd4168,15'd3848,15'd3528,15'd3208,15'd2888,15'd2568,15'd2248,15'd1928,15'd1608,15'd1288,15'd968,15'd648,15'd328,15'd8,
15'd25289,15'd24969,15'd24649,15'd24329,15'd24009,15'd23689,15'd23369,15'd23049,15'd22729,15'd22409,15'd22089,15'd21769,15'd21449,15'd21129,15'd20809,15'd20489,15'd20169,15'd19849,15'd19529,15'd19209,15'd18889,15'd18569,15'd18249,15'd17929,15'd17609,15'd17289,15'd16969,15'd16649,15'd16329,15'd16009,15'd15689,15'd15369,15'd15049,15'd14729,15'd14409,15'd14089,15'd13769,15'd13449,15'd13129,15'd12809,15'd12489,15'd12169,15'd11849,15'd11529,15'd11209,15'd10889,15'd10569,15'd10249,15'd9929,15'd9609,15'd9289,15'd8969,15'd8649,15'd8329,15'd8009,15'd7689,15'd7369,15'd7049,15'd6729,15'd6409,15'd6089,15'd5769,15'd5449,15'd5129,15'd4809,15'd4489,15'd4169,15'd3849,15'd3529,15'd3209,15'd2889,15'd2569,15'd2249,15'd1929,15'd1609,15'd1289,15'd969,15'd649,15'd329,15'd9,
15'd25290,15'd24970,15'd24650,15'd24330,15'd24010,15'd23690,15'd23370,15'd23050,15'd22730,15'd22410,15'd22090,15'd21770,15'd21450,15'd21130,15'd20810,15'd20490,15'd20170,15'd19850,15'd19530,15'd19210,15'd18890,15'd18570,15'd18250,15'd17930,15'd17610,15'd17290,15'd16970,15'd16650,15'd16330,15'd16010,15'd15690,15'd15370,15'd15050,15'd14730,15'd14410,15'd14090,15'd13770,15'd13450,15'd13130,15'd12810,15'd12490,15'd12170,15'd11850,15'd11530,15'd11210,15'd10890,15'd10570,15'd10250,15'd9930,15'd9610,15'd9290,15'd8970,15'd8650,15'd8330,15'd8010,15'd7690,15'd7370,15'd7050,15'd6730,15'd6410,15'd6090,15'd5770,15'd5450,15'd5130,15'd4810,15'd4490,15'd4170,15'd3850,15'd3530,15'd3210,15'd2890,15'd2570,15'd2250,15'd1930,15'd1610,15'd1290,15'd970,15'd650,15'd330,15'd10,
15'd25291,15'd24971,15'd24651,15'd24331,15'd24011,15'd23691,15'd23371,15'd23051,15'd22731,15'd22411,15'd22091,15'd21771,15'd21451,15'd21131,15'd20811,15'd20491,15'd20171,15'd19851,15'd19531,15'd19211,15'd18891,15'd18571,15'd18251,15'd17931,15'd17611,15'd17291,15'd16971,15'd16651,15'd16331,15'd16011,15'd15691,15'd15371,15'd15051,15'd14731,15'd14411,15'd14091,15'd13771,15'd13451,15'd13131,15'd12811,15'd12491,15'd12171,15'd11851,15'd11531,15'd11211,15'd10891,15'd10571,15'd10251,15'd9931,15'd9611,15'd9291,15'd8971,15'd8651,15'd8331,15'd8011,15'd7691,15'd7371,15'd7051,15'd6731,15'd6411,15'd6091,15'd5771,15'd5451,15'd5131,15'd4811,15'd4491,15'd4171,15'd3851,15'd3531,15'd3211,15'd2891,15'd2571,15'd2251,15'd1931,15'd1611,15'd1291,15'd971,15'd651,15'd331,15'd11,
15'd25292,15'd24972,15'd24652,15'd24332,15'd24012,15'd23692,15'd23372,15'd23052,15'd22732,15'd22412,15'd22092,15'd21772,15'd21452,15'd21132,15'd20812,15'd20492,15'd20172,15'd19852,15'd19532,15'd19212,15'd18892,15'd18572,15'd18252,15'd17932,15'd17612,15'd17292,15'd16972,15'd16652,15'd16332,15'd16012,15'd15692,15'd15372,15'd15052,15'd14732,15'd14412,15'd14092,15'd13772,15'd13452,15'd13132,15'd12812,15'd12492,15'd12172,15'd11852,15'd11532,15'd11212,15'd10892,15'd10572,15'd10252,15'd9932,15'd9612,15'd9292,15'd8972,15'd8652,15'd8332,15'd8012,15'd7692,15'd7372,15'd7052,15'd6732,15'd6412,15'd6092,15'd5772,15'd5452,15'd5132,15'd4812,15'd4492,15'd4172,15'd3852,15'd3532,15'd3212,15'd2892,15'd2572,15'd2252,15'd1932,15'd1612,15'd1292,15'd972,15'd652,15'd332,15'd12,
15'd25293,15'd24973,15'd24653,15'd24333,15'd24013,15'd23693,15'd23373,15'd23053,15'd22733,15'd22413,15'd22093,15'd21773,15'd21453,15'd21133,15'd20813,15'd20493,15'd20173,15'd19853,15'd19533,15'd19213,15'd18893,15'd18573,15'd18253,15'd17933,15'd17613,15'd17293,15'd16973,15'd16653,15'd16333,15'd16013,15'd15693,15'd15373,15'd15053,15'd14733,15'd14413,15'd14093,15'd13773,15'd13453,15'd13133,15'd12813,15'd12493,15'd12173,15'd11853,15'd11533,15'd11213,15'd10893,15'd10573,15'd10253,15'd9933,15'd9613,15'd9293,15'd8973,15'd8653,15'd8333,15'd8013,15'd7693,15'd7373,15'd7053,15'd6733,15'd6413,15'd6093,15'd5773,15'd5453,15'd5133,15'd4813,15'd4493,15'd4173,15'd3853,15'd3533,15'd3213,15'd2893,15'd2573,15'd2253,15'd1933,15'd1613,15'd1293,15'd973,15'd653,15'd333,15'd13,
15'd25294,15'd24974,15'd24654,15'd24334,15'd24014,15'd23694,15'd23374,15'd23054,15'd22734,15'd22414,15'd22094,15'd21774,15'd21454,15'd21134,15'd20814,15'd20494,15'd20174,15'd19854,15'd19534,15'd19214,15'd18894,15'd18574,15'd18254,15'd17934,15'd17614,15'd17294,15'd16974,15'd16654,15'd16334,15'd16014,15'd15694,15'd15374,15'd15054,15'd14734,15'd14414,15'd14094,15'd13774,15'd13454,15'd13134,15'd12814,15'd12494,15'd12174,15'd11854,15'd11534,15'd11214,15'd10894,15'd10574,15'd10254,15'd9934,15'd9614,15'd9294,15'd8974,15'd8654,15'd8334,15'd8014,15'd7694,15'd7374,15'd7054,15'd6734,15'd6414,15'd6094,15'd5774,15'd5454,15'd5134,15'd4814,15'd4494,15'd4174,15'd3854,15'd3534,15'd3214,15'd2894,15'd2574,15'd2254,15'd1934,15'd1614,15'd1294,15'd974,15'd654,15'd334,15'd14,
15'd25295,15'd24975,15'd24655,15'd24335,15'd24015,15'd23695,15'd23375,15'd23055,15'd22735,15'd22415,15'd22095,15'd21775,15'd21455,15'd21135,15'd20815,15'd20495,15'd20175,15'd19855,15'd19535,15'd19215,15'd18895,15'd18575,15'd18255,15'd17935,15'd17615,15'd17295,15'd16975,15'd16655,15'd16335,15'd16015,15'd15695,15'd15375,15'd15055,15'd14735,15'd14415,15'd14095,15'd13775,15'd13455,15'd13135,15'd12815,15'd12495,15'd12175,15'd11855,15'd11535,15'd11215,15'd10895,15'd10575,15'd10255,15'd9935,15'd9615,15'd9295,15'd8975,15'd8655,15'd8335,15'd8015,15'd7695,15'd7375,15'd7055,15'd6735,15'd6415,15'd6095,15'd5775,15'd5455,15'd5135,15'd4815,15'd4495,15'd4175,15'd3855,15'd3535,15'd3215,15'd2895,15'd2575,15'd2255,15'd1935,15'd1615,15'd1295,15'd975,15'd655,15'd335,15'd15,
15'd25296,15'd24976,15'd24656,15'd24336,15'd24016,15'd23696,15'd23376,15'd23056,15'd22736,15'd22416,15'd22096,15'd21776,15'd21456,15'd21136,15'd20816,15'd20496,15'd20176,15'd19856,15'd19536,15'd19216,15'd18896,15'd18576,15'd18256,15'd17936,15'd17616,15'd17296,15'd16976,15'd16656,15'd16336,15'd16016,15'd15696,15'd15376,15'd15056,15'd14736,15'd14416,15'd14096,15'd13776,15'd13456,15'd13136,15'd12816,15'd12496,15'd12176,15'd11856,15'd11536,15'd11216,15'd10896,15'd10576,15'd10256,15'd9936,15'd9616,15'd9296,15'd8976,15'd8656,15'd8336,15'd8016,15'd7696,15'd7376,15'd7056,15'd6736,15'd6416,15'd6096,15'd5776,15'd5456,15'd5136,15'd4816,15'd4496,15'd4176,15'd3856,15'd3536,15'd3216,15'd2896,15'd2576,15'd2256,15'd1936,15'd1616,15'd1296,15'd976,15'd656,15'd336,15'd16,
15'd25297,15'd24977,15'd24657,15'd24337,15'd24017,15'd23697,15'd23377,15'd23057,15'd22737,15'd22417,15'd22097,15'd21777,15'd21457,15'd21137,15'd20817,15'd20497,15'd20177,15'd19857,15'd19537,15'd19217,15'd18897,15'd18577,15'd18257,15'd17937,15'd17617,15'd17297,15'd16977,15'd16657,15'd16337,15'd16017,15'd15697,15'd15377,15'd15057,15'd14737,15'd14417,15'd14097,15'd13777,15'd13457,15'd13137,15'd12817,15'd12497,15'd12177,15'd11857,15'd11537,15'd11217,15'd10897,15'd10577,15'd10257,15'd9937,15'd9617,15'd9297,15'd8977,15'd8657,15'd8337,15'd8017,15'd7697,15'd7377,15'd7057,15'd6737,15'd6417,15'd6097,15'd5777,15'd5457,15'd5137,15'd4817,15'd4497,15'd4177,15'd3857,15'd3537,15'd3217,15'd2897,15'd2577,15'd2257,15'd1937,15'd1617,15'd1297,15'd977,15'd657,15'd337,15'd17,
15'd25298,15'd24978,15'd24658,15'd24338,15'd24018,15'd23698,15'd23378,15'd23058,15'd22738,15'd22418,15'd22098,15'd21778,15'd21458,15'd21138,15'd20818,15'd20498,15'd20178,15'd19858,15'd19538,15'd19218,15'd18898,15'd18578,15'd18258,15'd17938,15'd17618,15'd17298,15'd16978,15'd16658,15'd16338,15'd16018,15'd15698,15'd15378,15'd15058,15'd14738,15'd14418,15'd14098,15'd13778,15'd13458,15'd13138,15'd12818,15'd12498,15'd12178,15'd11858,15'd11538,15'd11218,15'd10898,15'd10578,15'd10258,15'd9938,15'd9618,15'd9298,15'd8978,15'd8658,15'd8338,15'd8018,15'd7698,15'd7378,15'd7058,15'd6738,15'd6418,15'd6098,15'd5778,15'd5458,15'd5138,15'd4818,15'd4498,15'd4178,15'd3858,15'd3538,15'd3218,15'd2898,15'd2578,15'd2258,15'd1938,15'd1618,15'd1298,15'd978,15'd658,15'd338,15'd18,
15'd25299,15'd24979,15'd24659,15'd24339,15'd24019,15'd23699,15'd23379,15'd23059,15'd22739,15'd22419,15'd22099,15'd21779,15'd21459,15'd21139,15'd20819,15'd20499,15'd20179,15'd19859,15'd19539,15'd19219,15'd18899,15'd18579,15'd18259,15'd17939,15'd17619,15'd17299,15'd16979,15'd16659,15'd16339,15'd16019,15'd15699,15'd15379,15'd15059,15'd14739,15'd14419,15'd14099,15'd13779,15'd13459,15'd13139,15'd12819,15'd12499,15'd12179,15'd11859,15'd11539,15'd11219,15'd10899,15'd10579,15'd10259,15'd9939,15'd9619,15'd9299,15'd8979,15'd8659,15'd8339,15'd8019,15'd7699,15'd7379,15'd7059,15'd6739,15'd6419,15'd6099,15'd5779,15'd5459,15'd5139,15'd4819,15'd4499,15'd4179,15'd3859,15'd3539,15'd3219,15'd2899,15'd2579,15'd2259,15'd1939,15'd1619,15'd1299,15'd979,15'd659,15'd339,15'd19,
15'd25300,15'd24980,15'd24660,15'd24340,15'd24020,15'd23700,15'd23380,15'd23060,15'd22740,15'd22420,15'd22100,15'd21780,15'd21460,15'd21140,15'd20820,15'd20500,15'd20180,15'd19860,15'd19540,15'd19220,15'd18900,15'd18580,15'd18260,15'd17940,15'd17620,15'd17300,15'd16980,15'd16660,15'd16340,15'd16020,15'd15700,15'd15380,15'd15060,15'd14740,15'd14420,15'd14100,15'd13780,15'd13460,15'd13140,15'd12820,15'd12500,15'd12180,15'd11860,15'd11540,15'd11220,15'd10900,15'd10580,15'd10260,15'd9940,15'd9620,15'd9300,15'd8980,15'd8660,15'd8340,15'd8020,15'd7700,15'd7380,15'd7060,15'd6740,15'd6420,15'd6100,15'd5780,15'd5460,15'd5140,15'd4820,15'd4500,15'd4180,15'd3860,15'd3540,15'd3220,15'd2900,15'd2580,15'd2260,15'd1940,15'd1620,15'd1300,15'd980,15'd660,15'd340,15'd20,
15'd25301,15'd24981,15'd24661,15'd24341,15'd24021,15'd23701,15'd23381,15'd23061,15'd22741,15'd22421,15'd22101,15'd21781,15'd21461,15'd21141,15'd20821,15'd20501,15'd20181,15'd19861,15'd19541,15'd19221,15'd18901,15'd18581,15'd18261,15'd17941,15'd17621,15'd17301,15'd16981,15'd16661,15'd16341,15'd16021,15'd15701,15'd15381,15'd15061,15'd14741,15'd14421,15'd14101,15'd13781,15'd13461,15'd13141,15'd12821,15'd12501,15'd12181,15'd11861,15'd11541,15'd11221,15'd10901,15'd10581,15'd10261,15'd9941,15'd9621,15'd9301,15'd8981,15'd8661,15'd8341,15'd8021,15'd7701,15'd7381,15'd7061,15'd6741,15'd6421,15'd6101,15'd5781,15'd5461,15'd5141,15'd4821,15'd4501,15'd4181,15'd3861,15'd3541,15'd3221,15'd2901,15'd2581,15'd2261,15'd1941,15'd1621,15'd1301,15'd981,15'd661,15'd341,15'd21,
15'd25302,15'd24982,15'd24662,15'd24342,15'd24022,15'd23702,15'd23382,15'd23062,15'd22742,15'd22422,15'd22102,15'd21782,15'd21462,15'd21142,15'd20822,15'd20502,15'd20182,15'd19862,15'd19542,15'd19222,15'd18902,15'd18582,15'd18262,15'd17942,15'd17622,15'd17302,15'd16982,15'd16662,15'd16342,15'd16022,15'd15702,15'd15382,15'd15062,15'd14742,15'd14422,15'd14102,15'd13782,15'd13462,15'd13142,15'd12822,15'd12502,15'd12182,15'd11862,15'd11542,15'd11222,15'd10902,15'd10582,15'd10262,15'd9942,15'd9622,15'd9302,15'd8982,15'd8662,15'd8342,15'd8022,15'd7702,15'd7382,15'd7062,15'd6742,15'd6422,15'd6102,15'd5782,15'd5462,15'd5142,15'd4822,15'd4502,15'd4182,15'd3862,15'd3542,15'd3222,15'd2902,15'd2582,15'd2262,15'd1942,15'd1622,15'd1302,15'd982,15'd662,15'd342,15'd22,
15'd25303,15'd24983,15'd24663,15'd24343,15'd24023,15'd23703,15'd23383,15'd23063,15'd22743,15'd22423,15'd22103,15'd21783,15'd21463,15'd21143,15'd20823,15'd20503,15'd20183,15'd19863,15'd19543,15'd19223,15'd18903,15'd18583,15'd18263,15'd17943,15'd17623,15'd17303,15'd16983,15'd16663,15'd16343,15'd16023,15'd15703,15'd15383,15'd15063,15'd14743,15'd14423,15'd14103,15'd13783,15'd13463,15'd13143,15'd12823,15'd12503,15'd12183,15'd11863,15'd11543,15'd11223,15'd10903,15'd10583,15'd10263,15'd9943,15'd9623,15'd9303,15'd8983,15'd8663,15'd8343,15'd8023,15'd7703,15'd7383,15'd7063,15'd6743,15'd6423,15'd6103,15'd5783,15'd5463,15'd5143,15'd4823,15'd4503,15'd4183,15'd3863,15'd3543,15'd3223,15'd2903,15'd2583,15'd2263,15'd1943,15'd1623,15'd1303,15'd983,15'd663,15'd343,15'd23,
15'd25304,15'd24984,15'd24664,15'd24344,15'd24024,15'd23704,15'd23384,15'd23064,15'd22744,15'd22424,15'd22104,15'd21784,15'd21464,15'd21144,15'd20824,15'd20504,15'd20184,15'd19864,15'd19544,15'd19224,15'd18904,15'd18584,15'd18264,15'd17944,15'd17624,15'd17304,15'd16984,15'd16664,15'd16344,15'd16024,15'd15704,15'd15384,15'd15064,15'd14744,15'd14424,15'd14104,15'd13784,15'd13464,15'd13144,15'd12824,15'd12504,15'd12184,15'd11864,15'd11544,15'd11224,15'd10904,15'd10584,15'd10264,15'd9944,15'd9624,15'd9304,15'd8984,15'd8664,15'd8344,15'd8024,15'd7704,15'd7384,15'd7064,15'd6744,15'd6424,15'd6104,15'd5784,15'd5464,15'd5144,15'd4824,15'd4504,15'd4184,15'd3864,15'd3544,15'd3224,15'd2904,15'd2584,15'd2264,15'd1944,15'd1624,15'd1304,15'd984,15'd664,15'd344,15'd24,
15'd25305,15'd24985,15'd24665,15'd24345,15'd24025,15'd23705,15'd23385,15'd23065,15'd22745,15'd22425,15'd22105,15'd21785,15'd21465,15'd21145,15'd20825,15'd20505,15'd20185,15'd19865,15'd19545,15'd19225,15'd18905,15'd18585,15'd18265,15'd17945,15'd17625,15'd17305,15'd16985,15'd16665,15'd16345,15'd16025,15'd15705,15'd15385,15'd15065,15'd14745,15'd14425,15'd14105,15'd13785,15'd13465,15'd13145,15'd12825,15'd12505,15'd12185,15'd11865,15'd11545,15'd11225,15'd10905,15'd10585,15'd10265,15'd9945,15'd9625,15'd9305,15'd8985,15'd8665,15'd8345,15'd8025,15'd7705,15'd7385,15'd7065,15'd6745,15'd6425,15'd6105,15'd5785,15'd5465,15'd5145,15'd4825,15'd4505,15'd4185,15'd3865,15'd3545,15'd3225,15'd2905,15'd2585,15'd2265,15'd1945,15'd1625,15'd1305,15'd985,15'd665,15'd345,15'd25,
15'd25306,15'd24986,15'd24666,15'd24346,15'd24026,15'd23706,15'd23386,15'd23066,15'd22746,15'd22426,15'd22106,15'd21786,15'd21466,15'd21146,15'd20826,15'd20506,15'd20186,15'd19866,15'd19546,15'd19226,15'd18906,15'd18586,15'd18266,15'd17946,15'd17626,15'd17306,15'd16986,15'd16666,15'd16346,15'd16026,15'd15706,15'd15386,15'd15066,15'd14746,15'd14426,15'd14106,15'd13786,15'd13466,15'd13146,15'd12826,15'd12506,15'd12186,15'd11866,15'd11546,15'd11226,15'd10906,15'd10586,15'd10266,15'd9946,15'd9626,15'd9306,15'd8986,15'd8666,15'd8346,15'd8026,15'd7706,15'd7386,15'd7066,15'd6746,15'd6426,15'd6106,15'd5786,15'd5466,15'd5146,15'd4826,15'd4506,15'd4186,15'd3866,15'd3546,15'd3226,15'd2906,15'd2586,15'd2266,15'd1946,15'd1626,15'd1306,15'd986,15'd666,15'd346,15'd26,
15'd25307,15'd24987,15'd24667,15'd24347,15'd24027,15'd23707,15'd23387,15'd23067,15'd22747,15'd22427,15'd22107,15'd21787,15'd21467,15'd21147,15'd20827,15'd20507,15'd20187,15'd19867,15'd19547,15'd19227,15'd18907,15'd18587,15'd18267,15'd17947,15'd17627,15'd17307,15'd16987,15'd16667,15'd16347,15'd16027,15'd15707,15'd15387,15'd15067,15'd14747,15'd14427,15'd14107,15'd13787,15'd13467,15'd13147,15'd12827,15'd12507,15'd12187,15'd11867,15'd11547,15'd11227,15'd10907,15'd10587,15'd10267,15'd9947,15'd9627,15'd9307,15'd8987,15'd8667,15'd8347,15'd8027,15'd7707,15'd7387,15'd7067,15'd6747,15'd6427,15'd6107,15'd5787,15'd5467,15'd5147,15'd4827,15'd4507,15'd4187,15'd3867,15'd3547,15'd3227,15'd2907,15'd2587,15'd2267,15'd1947,15'd1627,15'd1307,15'd987,15'd667,15'd347,15'd27,
15'd25308,15'd24988,15'd24668,15'd24348,15'd24028,15'd23708,15'd23388,15'd23068,15'd22748,15'd22428,15'd22108,15'd21788,15'd21468,15'd21148,15'd20828,15'd20508,15'd20188,15'd19868,15'd19548,15'd19228,15'd18908,15'd18588,15'd18268,15'd17948,15'd17628,15'd17308,15'd16988,15'd16668,15'd16348,15'd16028,15'd15708,15'd15388,15'd15068,15'd14748,15'd14428,15'd14108,15'd13788,15'd13468,15'd13148,15'd12828,15'd12508,15'd12188,15'd11868,15'd11548,15'd11228,15'd10908,15'd10588,15'd10268,15'd9948,15'd9628,15'd9308,15'd8988,15'd8668,15'd8348,15'd8028,15'd7708,15'd7388,15'd7068,15'd6748,15'd6428,15'd6108,15'd5788,15'd5468,15'd5148,15'd4828,15'd4508,15'd4188,15'd3868,15'd3548,15'd3228,15'd2908,15'd2588,15'd2268,15'd1948,15'd1628,15'd1308,15'd988,15'd668,15'd348,15'd28,
15'd25309,15'd24989,15'd24669,15'd24349,15'd24029,15'd23709,15'd23389,15'd23069,15'd22749,15'd22429,15'd22109,15'd21789,15'd21469,15'd21149,15'd20829,15'd20509,15'd20189,15'd19869,15'd19549,15'd19229,15'd18909,15'd18589,15'd18269,15'd17949,15'd17629,15'd17309,15'd16989,15'd16669,15'd16349,15'd16029,15'd15709,15'd15389,15'd15069,15'd14749,15'd14429,15'd14109,15'd13789,15'd13469,15'd13149,15'd12829,15'd12509,15'd12189,15'd11869,15'd11549,15'd11229,15'd10909,15'd10589,15'd10269,15'd9949,15'd9629,15'd9309,15'd8989,15'd8669,15'd8349,15'd8029,15'd7709,15'd7389,15'd7069,15'd6749,15'd6429,15'd6109,15'd5789,15'd5469,15'd5149,15'd4829,15'd4509,15'd4189,15'd3869,15'd3549,15'd3229,15'd2909,15'd2589,15'd2269,15'd1949,15'd1629,15'd1309,15'd989,15'd669,15'd349,15'd29,
15'd25310,15'd24990,15'd24670,15'd24350,15'd24030,15'd23710,15'd23390,15'd23070,15'd22750,15'd22430,15'd22110,15'd21790,15'd21470,15'd21150,15'd20830,15'd20510,15'd20190,15'd19870,15'd19550,15'd19230,15'd18910,15'd18590,15'd18270,15'd17950,15'd17630,15'd17310,15'd16990,15'd16670,15'd16350,15'd16030,15'd15710,15'd15390,15'd15070,15'd14750,15'd14430,15'd14110,15'd13790,15'd13470,15'd13150,15'd12830,15'd12510,15'd12190,15'd11870,15'd11550,15'd11230,15'd10910,15'd10590,15'd10270,15'd9950,15'd9630,15'd9310,15'd8990,15'd8670,15'd8350,15'd8030,15'd7710,15'd7390,15'd7070,15'd6750,15'd6430,15'd6110,15'd5790,15'd5470,15'd5150,15'd4830,15'd4510,15'd4190,15'd3870,15'd3550,15'd3230,15'd2910,15'd2590,15'd2270,15'd1950,15'd1630,15'd1310,15'd990,15'd670,15'd350,15'd30,
15'd25311,15'd24991,15'd24671,15'd24351,15'd24031,15'd23711,15'd23391,15'd23071,15'd22751,15'd22431,15'd22111,15'd21791,15'd21471,15'd21151,15'd20831,15'd20511,15'd20191,15'd19871,15'd19551,15'd19231,15'd18911,15'd18591,15'd18271,15'd17951,15'd17631,15'd17311,15'd16991,15'd16671,15'd16351,15'd16031,15'd15711,15'd15391,15'd15071,15'd14751,15'd14431,15'd14111,15'd13791,15'd13471,15'd13151,15'd12831,15'd12511,15'd12191,15'd11871,15'd11551,15'd11231,15'd10911,15'd10591,15'd10271,15'd9951,15'd9631,15'd9311,15'd8991,15'd8671,15'd8351,15'd8031,15'd7711,15'd7391,15'd7071,15'd6751,15'd6431,15'd6111,15'd5791,15'd5471,15'd5151,15'd4831,15'd4511,15'd4191,15'd3871,15'd3551,15'd3231,15'd2911,15'd2591,15'd2271,15'd1951,15'd1631,15'd1311,15'd991,15'd671,15'd351,15'd31,
15'd25312,15'd24992,15'd24672,15'd24352,15'd24032,15'd23712,15'd23392,15'd23072,15'd22752,15'd22432,15'd22112,15'd21792,15'd21472,15'd21152,15'd20832,15'd20512,15'd20192,15'd19872,15'd19552,15'd19232,15'd18912,15'd18592,15'd18272,15'd17952,15'd17632,15'd17312,15'd16992,15'd16672,15'd16352,15'd16032,15'd15712,15'd15392,15'd15072,15'd14752,15'd14432,15'd14112,15'd13792,15'd13472,15'd13152,15'd12832,15'd12512,15'd12192,15'd11872,15'd11552,15'd11232,15'd10912,15'd10592,15'd10272,15'd9952,15'd9632,15'd9312,15'd8992,15'd8672,15'd8352,15'd8032,15'd7712,15'd7392,15'd7072,15'd6752,15'd6432,15'd6112,15'd5792,15'd5472,15'd5152,15'd4832,15'd4512,15'd4192,15'd3872,15'd3552,15'd3232,15'd2912,15'd2592,15'd2272,15'd1952,15'd1632,15'd1312,15'd992,15'd672,15'd352,15'd32,
15'd25313,15'd24993,15'd24673,15'd24353,15'd24033,15'd23713,15'd23393,15'd23073,15'd22753,15'd22433,15'd22113,15'd21793,15'd21473,15'd21153,15'd20833,15'd20513,15'd20193,15'd19873,15'd19553,15'd19233,15'd18913,15'd18593,15'd18273,15'd17953,15'd17633,15'd17313,15'd16993,15'd16673,15'd16353,15'd16033,15'd15713,15'd15393,15'd15073,15'd14753,15'd14433,15'd14113,15'd13793,15'd13473,15'd13153,15'd12833,15'd12513,15'd12193,15'd11873,15'd11553,15'd11233,15'd10913,15'd10593,15'd10273,15'd9953,15'd9633,15'd9313,15'd8993,15'd8673,15'd8353,15'd8033,15'd7713,15'd7393,15'd7073,15'd6753,15'd6433,15'd6113,15'd5793,15'd5473,15'd5153,15'd4833,15'd4513,15'd4193,15'd3873,15'd3553,15'd3233,15'd2913,15'd2593,15'd2273,15'd1953,15'd1633,15'd1313,15'd993,15'd673,15'd353,15'd33,
15'd25314,15'd24994,15'd24674,15'd24354,15'd24034,15'd23714,15'd23394,15'd23074,15'd22754,15'd22434,15'd22114,15'd21794,15'd21474,15'd21154,15'd20834,15'd20514,15'd20194,15'd19874,15'd19554,15'd19234,15'd18914,15'd18594,15'd18274,15'd17954,15'd17634,15'd17314,15'd16994,15'd16674,15'd16354,15'd16034,15'd15714,15'd15394,15'd15074,15'd14754,15'd14434,15'd14114,15'd13794,15'd13474,15'd13154,15'd12834,15'd12514,15'd12194,15'd11874,15'd11554,15'd11234,15'd10914,15'd10594,15'd10274,15'd9954,15'd9634,15'd9314,15'd8994,15'd8674,15'd8354,15'd8034,15'd7714,15'd7394,15'd7074,15'd6754,15'd6434,15'd6114,15'd5794,15'd5474,15'd5154,15'd4834,15'd4514,15'd4194,15'd3874,15'd3554,15'd3234,15'd2914,15'd2594,15'd2274,15'd1954,15'd1634,15'd1314,15'd994,15'd674,15'd354,15'd34,
15'd25315,15'd24995,15'd24675,15'd24355,15'd24035,15'd23715,15'd23395,15'd23075,15'd22755,15'd22435,15'd22115,15'd21795,15'd21475,15'd21155,15'd20835,15'd20515,15'd20195,15'd19875,15'd19555,15'd19235,15'd18915,15'd18595,15'd18275,15'd17955,15'd17635,15'd17315,15'd16995,15'd16675,15'd16355,15'd16035,15'd15715,15'd15395,15'd15075,15'd14755,15'd14435,15'd14115,15'd13795,15'd13475,15'd13155,15'd12835,15'd12515,15'd12195,15'd11875,15'd11555,15'd11235,15'd10915,15'd10595,15'd10275,15'd9955,15'd9635,15'd9315,15'd8995,15'd8675,15'd8355,15'd8035,15'd7715,15'd7395,15'd7075,15'd6755,15'd6435,15'd6115,15'd5795,15'd5475,15'd5155,15'd4835,15'd4515,15'd4195,15'd3875,15'd3555,15'd3235,15'd2915,15'd2595,15'd2275,15'd1955,15'd1635,15'd1315,15'd995,15'd675,15'd355,15'd35,
15'd25316,15'd24996,15'd24676,15'd24356,15'd24036,15'd23716,15'd23396,15'd23076,15'd22756,15'd22436,15'd22116,15'd21796,15'd21476,15'd21156,15'd20836,15'd20516,15'd20196,15'd19876,15'd19556,15'd19236,15'd18916,15'd18596,15'd18276,15'd17956,15'd17636,15'd17316,15'd16996,15'd16676,15'd16356,15'd16036,15'd15716,15'd15396,15'd15076,15'd14756,15'd14436,15'd14116,15'd13796,15'd13476,15'd13156,15'd12836,15'd12516,15'd12196,15'd11876,15'd11556,15'd11236,15'd10916,15'd10596,15'd10276,15'd9956,15'd9636,15'd9316,15'd8996,15'd8676,15'd8356,15'd8036,15'd7716,15'd7396,15'd7076,15'd6756,15'd6436,15'd6116,15'd5796,15'd5476,15'd5156,15'd4836,15'd4516,15'd4196,15'd3876,15'd3556,15'd3236,15'd2916,15'd2596,15'd2276,15'd1956,15'd1636,15'd1316,15'd996,15'd676,15'd356,15'd36,
15'd25317,15'd24997,15'd24677,15'd24357,15'd24037,15'd23717,15'd23397,15'd23077,15'd22757,15'd22437,15'd22117,15'd21797,15'd21477,15'd21157,15'd20837,15'd20517,15'd20197,15'd19877,15'd19557,15'd19237,15'd18917,15'd18597,15'd18277,15'd17957,15'd17637,15'd17317,15'd16997,15'd16677,15'd16357,15'd16037,15'd15717,15'd15397,15'd15077,15'd14757,15'd14437,15'd14117,15'd13797,15'd13477,15'd13157,15'd12837,15'd12517,15'd12197,15'd11877,15'd11557,15'd11237,15'd10917,15'd10597,15'd10277,15'd9957,15'd9637,15'd9317,15'd8997,15'd8677,15'd8357,15'd8037,15'd7717,15'd7397,15'd7077,15'd6757,15'd6437,15'd6117,15'd5797,15'd5477,15'd5157,15'd4837,15'd4517,15'd4197,15'd3877,15'd3557,15'd3237,15'd2917,15'd2597,15'd2277,15'd1957,15'd1637,15'd1317,15'd997,15'd677,15'd357,15'd37,
15'd25318,15'd24998,15'd24678,15'd24358,15'd24038,15'd23718,15'd23398,15'd23078,15'd22758,15'd22438,15'd22118,15'd21798,15'd21478,15'd21158,15'd20838,15'd20518,15'd20198,15'd19878,15'd19558,15'd19238,15'd18918,15'd18598,15'd18278,15'd17958,15'd17638,15'd17318,15'd16998,15'd16678,15'd16358,15'd16038,15'd15718,15'd15398,15'd15078,15'd14758,15'd14438,15'd14118,15'd13798,15'd13478,15'd13158,15'd12838,15'd12518,15'd12198,15'd11878,15'd11558,15'd11238,15'd10918,15'd10598,15'd10278,15'd9958,15'd9638,15'd9318,15'd8998,15'd8678,15'd8358,15'd8038,15'd7718,15'd7398,15'd7078,15'd6758,15'd6438,15'd6118,15'd5798,15'd5478,15'd5158,15'd4838,15'd4518,15'd4198,15'd3878,15'd3558,15'd3238,15'd2918,15'd2598,15'd2278,15'd1958,15'd1638,15'd1318,15'd998,15'd678,15'd358,15'd38,
15'd25319,15'd24999,15'd24679,15'd24359,15'd24039,15'd23719,15'd23399,15'd23079,15'd22759,15'd22439,15'd22119,15'd21799,15'd21479,15'd21159,15'd20839,15'd20519,15'd20199,15'd19879,15'd19559,15'd19239,15'd18919,15'd18599,15'd18279,15'd17959,15'd17639,15'd17319,15'd16999,15'd16679,15'd16359,15'd16039,15'd15719,15'd15399,15'd15079,15'd14759,15'd14439,15'd14119,15'd13799,15'd13479,15'd13159,15'd12839,15'd12519,15'd12199,15'd11879,15'd11559,15'd11239,15'd10919,15'd10599,15'd10279,15'd9959,15'd9639,15'd9319,15'd8999,15'd8679,15'd8359,15'd8039,15'd7719,15'd7399,15'd7079,15'd6759,15'd6439,15'd6119,15'd5799,15'd5479,15'd5159,15'd4839,15'd4519,15'd4199,15'd3879,15'd3559,15'd3239,15'd2919,15'd2599,15'd2279,15'd1959,15'd1639,15'd1319,15'd999,15'd679,15'd359,15'd39,
15'd25320,15'd25000,15'd24680,15'd24360,15'd24040,15'd23720,15'd23400,15'd23080,15'd22760,15'd22440,15'd22120,15'd21800,15'd21480,15'd21160,15'd20840,15'd20520,15'd20200,15'd19880,15'd19560,15'd19240,15'd18920,15'd18600,15'd18280,15'd17960,15'd17640,15'd17320,15'd17000,15'd16680,15'd16360,15'd16040,15'd15720,15'd15400,15'd15080,15'd14760,15'd14440,15'd14120,15'd13800,15'd13480,15'd13160,15'd12840,15'd12520,15'd12200,15'd11880,15'd11560,15'd11240,15'd10920,15'd10600,15'd10280,15'd9960,15'd9640,15'd9320,15'd9000,15'd8680,15'd8360,15'd8040,15'd7720,15'd7400,15'd7080,15'd6760,15'd6440,15'd6120,15'd5800,15'd5480,15'd5160,15'd4840,15'd4520,15'd4200,15'd3880,15'd3560,15'd3240,15'd2920,15'd2600,15'd2280,15'd1960,15'd1640,15'd1320,15'd1000,15'd680,15'd360,15'd40,
15'd25321,15'd25001,15'd24681,15'd24361,15'd24041,15'd23721,15'd23401,15'd23081,15'd22761,15'd22441,15'd22121,15'd21801,15'd21481,15'd21161,15'd20841,15'd20521,15'd20201,15'd19881,15'd19561,15'd19241,15'd18921,15'd18601,15'd18281,15'd17961,15'd17641,15'd17321,15'd17001,15'd16681,15'd16361,15'd16041,15'd15721,15'd15401,15'd15081,15'd14761,15'd14441,15'd14121,15'd13801,15'd13481,15'd13161,15'd12841,15'd12521,15'd12201,15'd11881,15'd11561,15'd11241,15'd10921,15'd10601,15'd10281,15'd9961,15'd9641,15'd9321,15'd9001,15'd8681,15'd8361,15'd8041,15'd7721,15'd7401,15'd7081,15'd6761,15'd6441,15'd6121,15'd5801,15'd5481,15'd5161,15'd4841,15'd4521,15'd4201,15'd3881,15'd3561,15'd3241,15'd2921,15'd2601,15'd2281,15'd1961,15'd1641,15'd1321,15'd1001,15'd681,15'd361,15'd41,
15'd25322,15'd25002,15'd24682,15'd24362,15'd24042,15'd23722,15'd23402,15'd23082,15'd22762,15'd22442,15'd22122,15'd21802,15'd21482,15'd21162,15'd20842,15'd20522,15'd20202,15'd19882,15'd19562,15'd19242,15'd18922,15'd18602,15'd18282,15'd17962,15'd17642,15'd17322,15'd17002,15'd16682,15'd16362,15'd16042,15'd15722,15'd15402,15'd15082,15'd14762,15'd14442,15'd14122,15'd13802,15'd13482,15'd13162,15'd12842,15'd12522,15'd12202,15'd11882,15'd11562,15'd11242,15'd10922,15'd10602,15'd10282,15'd9962,15'd9642,15'd9322,15'd9002,15'd8682,15'd8362,15'd8042,15'd7722,15'd7402,15'd7082,15'd6762,15'd6442,15'd6122,15'd5802,15'd5482,15'd5162,15'd4842,15'd4522,15'd4202,15'd3882,15'd3562,15'd3242,15'd2922,15'd2602,15'd2282,15'd1962,15'd1642,15'd1322,15'd1002,15'd682,15'd362,15'd42,
15'd25323,15'd25003,15'd24683,15'd24363,15'd24043,15'd23723,15'd23403,15'd23083,15'd22763,15'd22443,15'd22123,15'd21803,15'd21483,15'd21163,15'd20843,15'd20523,15'd20203,15'd19883,15'd19563,15'd19243,15'd18923,15'd18603,15'd18283,15'd17963,15'd17643,15'd17323,15'd17003,15'd16683,15'd16363,15'd16043,15'd15723,15'd15403,15'd15083,15'd14763,15'd14443,15'd14123,15'd13803,15'd13483,15'd13163,15'd12843,15'd12523,15'd12203,15'd11883,15'd11563,15'd11243,15'd10923,15'd10603,15'd10283,15'd9963,15'd9643,15'd9323,15'd9003,15'd8683,15'd8363,15'd8043,15'd7723,15'd7403,15'd7083,15'd6763,15'd6443,15'd6123,15'd5803,15'd5483,15'd5163,15'd4843,15'd4523,15'd4203,15'd3883,15'd3563,15'd3243,15'd2923,15'd2603,15'd2283,15'd1963,15'd1643,15'd1323,15'd1003,15'd683,15'd363,15'd43,
15'd25324,15'd25004,15'd24684,15'd24364,15'd24044,15'd23724,15'd23404,15'd23084,15'd22764,15'd22444,15'd22124,15'd21804,15'd21484,15'd21164,15'd20844,15'd20524,15'd20204,15'd19884,15'd19564,15'd19244,15'd18924,15'd18604,15'd18284,15'd17964,15'd17644,15'd17324,15'd17004,15'd16684,15'd16364,15'd16044,15'd15724,15'd15404,15'd15084,15'd14764,15'd14444,15'd14124,15'd13804,15'd13484,15'd13164,15'd12844,15'd12524,15'd12204,15'd11884,15'd11564,15'd11244,15'd10924,15'd10604,15'd10284,15'd9964,15'd9644,15'd9324,15'd9004,15'd8684,15'd8364,15'd8044,15'd7724,15'd7404,15'd7084,15'd6764,15'd6444,15'd6124,15'd5804,15'd5484,15'd5164,15'd4844,15'd4524,15'd4204,15'd3884,15'd3564,15'd3244,15'd2924,15'd2604,15'd2284,15'd1964,15'd1644,15'd1324,15'd1004,15'd684,15'd364,15'd44,
15'd25325,15'd25005,15'd24685,15'd24365,15'd24045,15'd23725,15'd23405,15'd23085,15'd22765,15'd22445,15'd22125,15'd21805,15'd21485,15'd21165,15'd20845,15'd20525,15'd20205,15'd19885,15'd19565,15'd19245,15'd18925,15'd18605,15'd18285,15'd17965,15'd17645,15'd17325,15'd17005,15'd16685,15'd16365,15'd16045,15'd15725,15'd15405,15'd15085,15'd14765,15'd14445,15'd14125,15'd13805,15'd13485,15'd13165,15'd12845,15'd12525,15'd12205,15'd11885,15'd11565,15'd11245,15'd10925,15'd10605,15'd10285,15'd9965,15'd9645,15'd9325,15'd9005,15'd8685,15'd8365,15'd8045,15'd7725,15'd7405,15'd7085,15'd6765,15'd6445,15'd6125,15'd5805,15'd5485,15'd5165,15'd4845,15'd4525,15'd4205,15'd3885,15'd3565,15'd3245,15'd2925,15'd2605,15'd2285,15'd1965,15'd1645,15'd1325,15'd1005,15'd685,15'd365,15'd45,
15'd25326,15'd25006,15'd24686,15'd24366,15'd24046,15'd23726,15'd23406,15'd23086,15'd22766,15'd22446,15'd22126,15'd21806,15'd21486,15'd21166,15'd20846,15'd20526,15'd20206,15'd19886,15'd19566,15'd19246,15'd18926,15'd18606,15'd18286,15'd17966,15'd17646,15'd17326,15'd17006,15'd16686,15'd16366,15'd16046,15'd15726,15'd15406,15'd15086,15'd14766,15'd14446,15'd14126,15'd13806,15'd13486,15'd13166,15'd12846,15'd12526,15'd12206,15'd11886,15'd11566,15'd11246,15'd10926,15'd10606,15'd10286,15'd9966,15'd9646,15'd9326,15'd9006,15'd8686,15'd8366,15'd8046,15'd7726,15'd7406,15'd7086,15'd6766,15'd6446,15'd6126,15'd5806,15'd5486,15'd5166,15'd4846,15'd4526,15'd4206,15'd3886,15'd3566,15'd3246,15'd2926,15'd2606,15'd2286,15'd1966,15'd1646,15'd1326,15'd1006,15'd686,15'd366,15'd46,
15'd25327,15'd25007,15'd24687,15'd24367,15'd24047,15'd23727,15'd23407,15'd23087,15'd22767,15'd22447,15'd22127,15'd21807,15'd21487,15'd21167,15'd20847,15'd20527,15'd20207,15'd19887,15'd19567,15'd19247,15'd18927,15'd18607,15'd18287,15'd17967,15'd17647,15'd17327,15'd17007,15'd16687,15'd16367,15'd16047,15'd15727,15'd15407,15'd15087,15'd14767,15'd14447,15'd14127,15'd13807,15'd13487,15'd13167,15'd12847,15'd12527,15'd12207,15'd11887,15'd11567,15'd11247,15'd10927,15'd10607,15'd10287,15'd9967,15'd9647,15'd9327,15'd9007,15'd8687,15'd8367,15'd8047,15'd7727,15'd7407,15'd7087,15'd6767,15'd6447,15'd6127,15'd5807,15'd5487,15'd5167,15'd4847,15'd4527,15'd4207,15'd3887,15'd3567,15'd3247,15'd2927,15'd2607,15'd2287,15'd1967,15'd1647,15'd1327,15'd1007,15'd687,15'd367,15'd47,
15'd25328,15'd25008,15'd24688,15'd24368,15'd24048,15'd23728,15'd23408,15'd23088,15'd22768,15'd22448,15'd22128,15'd21808,15'd21488,15'd21168,15'd20848,15'd20528,15'd20208,15'd19888,15'd19568,15'd19248,15'd18928,15'd18608,15'd18288,15'd17968,15'd17648,15'd17328,15'd17008,15'd16688,15'd16368,15'd16048,15'd15728,15'd15408,15'd15088,15'd14768,15'd14448,15'd14128,15'd13808,15'd13488,15'd13168,15'd12848,15'd12528,15'd12208,15'd11888,15'd11568,15'd11248,15'd10928,15'd10608,15'd10288,15'd9968,15'd9648,15'd9328,15'd9008,15'd8688,15'd8368,15'd8048,15'd7728,15'd7408,15'd7088,15'd6768,15'd6448,15'd6128,15'd5808,15'd5488,15'd5168,15'd4848,15'd4528,15'd4208,15'd3888,15'd3568,15'd3248,15'd2928,15'd2608,15'd2288,15'd1968,15'd1648,15'd1328,15'd1008,15'd688,15'd368,15'd48,
15'd25329,15'd25009,15'd24689,15'd24369,15'd24049,15'd23729,15'd23409,15'd23089,15'd22769,15'd22449,15'd22129,15'd21809,15'd21489,15'd21169,15'd20849,15'd20529,15'd20209,15'd19889,15'd19569,15'd19249,15'd18929,15'd18609,15'd18289,15'd17969,15'd17649,15'd17329,15'd17009,15'd16689,15'd16369,15'd16049,15'd15729,15'd15409,15'd15089,15'd14769,15'd14449,15'd14129,15'd13809,15'd13489,15'd13169,15'd12849,15'd12529,15'd12209,15'd11889,15'd11569,15'd11249,15'd10929,15'd10609,15'd10289,15'd9969,15'd9649,15'd9329,15'd9009,15'd8689,15'd8369,15'd8049,15'd7729,15'd7409,15'd7089,15'd6769,15'd6449,15'd6129,15'd5809,15'd5489,15'd5169,15'd4849,15'd4529,15'd4209,15'd3889,15'd3569,15'd3249,15'd2929,15'd2609,15'd2289,15'd1969,15'd1649,15'd1329,15'd1009,15'd689,15'd369,15'd49,
15'd25330,15'd25010,15'd24690,15'd24370,15'd24050,15'd23730,15'd23410,15'd23090,15'd22770,15'd22450,15'd22130,15'd21810,15'd21490,15'd21170,15'd20850,15'd20530,15'd20210,15'd19890,15'd19570,15'd19250,15'd18930,15'd18610,15'd18290,15'd17970,15'd17650,15'd17330,15'd17010,15'd16690,15'd16370,15'd16050,15'd15730,15'd15410,15'd15090,15'd14770,15'd14450,15'd14130,15'd13810,15'd13490,15'd13170,15'd12850,15'd12530,15'd12210,15'd11890,15'd11570,15'd11250,15'd10930,15'd10610,15'd10290,15'd9970,15'd9650,15'd9330,15'd9010,15'd8690,15'd8370,15'd8050,15'd7730,15'd7410,15'd7090,15'd6770,15'd6450,15'd6130,15'd5810,15'd5490,15'd5170,15'd4850,15'd4530,15'd4210,15'd3890,15'd3570,15'd3250,15'd2930,15'd2610,15'd2290,15'd1970,15'd1650,15'd1330,15'd1010,15'd690,15'd370,15'd50,
15'd25331,15'd25011,15'd24691,15'd24371,15'd24051,15'd23731,15'd23411,15'd23091,15'd22771,15'd22451,15'd22131,15'd21811,15'd21491,15'd21171,15'd20851,15'd20531,15'd20211,15'd19891,15'd19571,15'd19251,15'd18931,15'd18611,15'd18291,15'd17971,15'd17651,15'd17331,15'd17011,15'd16691,15'd16371,15'd16051,15'd15731,15'd15411,15'd15091,15'd14771,15'd14451,15'd14131,15'd13811,15'd13491,15'd13171,15'd12851,15'd12531,15'd12211,15'd11891,15'd11571,15'd11251,15'd10931,15'd10611,15'd10291,15'd9971,15'd9651,15'd9331,15'd9011,15'd8691,15'd8371,15'd8051,15'd7731,15'd7411,15'd7091,15'd6771,15'd6451,15'd6131,15'd5811,15'd5491,15'd5171,15'd4851,15'd4531,15'd4211,15'd3891,15'd3571,15'd3251,15'd2931,15'd2611,15'd2291,15'd1971,15'd1651,15'd1331,15'd1011,15'd691,15'd371,15'd51,
15'd25332,15'd25012,15'd24692,15'd24372,15'd24052,15'd23732,15'd23412,15'd23092,15'd22772,15'd22452,15'd22132,15'd21812,15'd21492,15'd21172,15'd20852,15'd20532,15'd20212,15'd19892,15'd19572,15'd19252,15'd18932,15'd18612,15'd18292,15'd17972,15'd17652,15'd17332,15'd17012,15'd16692,15'd16372,15'd16052,15'd15732,15'd15412,15'd15092,15'd14772,15'd14452,15'd14132,15'd13812,15'd13492,15'd13172,15'd12852,15'd12532,15'd12212,15'd11892,15'd11572,15'd11252,15'd10932,15'd10612,15'd10292,15'd9972,15'd9652,15'd9332,15'd9012,15'd8692,15'd8372,15'd8052,15'd7732,15'd7412,15'd7092,15'd6772,15'd6452,15'd6132,15'd5812,15'd5492,15'd5172,15'd4852,15'd4532,15'd4212,15'd3892,15'd3572,15'd3252,15'd2932,15'd2612,15'd2292,15'd1972,15'd1652,15'd1332,15'd1012,15'd692,15'd372,15'd52,
15'd25333,15'd25013,15'd24693,15'd24373,15'd24053,15'd23733,15'd23413,15'd23093,15'd22773,15'd22453,15'd22133,15'd21813,15'd21493,15'd21173,15'd20853,15'd20533,15'd20213,15'd19893,15'd19573,15'd19253,15'd18933,15'd18613,15'd18293,15'd17973,15'd17653,15'd17333,15'd17013,15'd16693,15'd16373,15'd16053,15'd15733,15'd15413,15'd15093,15'd14773,15'd14453,15'd14133,15'd13813,15'd13493,15'd13173,15'd12853,15'd12533,15'd12213,15'd11893,15'd11573,15'd11253,15'd10933,15'd10613,15'd10293,15'd9973,15'd9653,15'd9333,15'd9013,15'd8693,15'd8373,15'd8053,15'd7733,15'd7413,15'd7093,15'd6773,15'd6453,15'd6133,15'd5813,15'd5493,15'd5173,15'd4853,15'd4533,15'd4213,15'd3893,15'd3573,15'd3253,15'd2933,15'd2613,15'd2293,15'd1973,15'd1653,15'd1333,15'd1013,15'd693,15'd373,15'd53,
15'd25334,15'd25014,15'd24694,15'd24374,15'd24054,15'd23734,15'd23414,15'd23094,15'd22774,15'd22454,15'd22134,15'd21814,15'd21494,15'd21174,15'd20854,15'd20534,15'd20214,15'd19894,15'd19574,15'd19254,15'd18934,15'd18614,15'd18294,15'd17974,15'd17654,15'd17334,15'd17014,15'd16694,15'd16374,15'd16054,15'd15734,15'd15414,15'd15094,15'd14774,15'd14454,15'd14134,15'd13814,15'd13494,15'd13174,15'd12854,15'd12534,15'd12214,15'd11894,15'd11574,15'd11254,15'd10934,15'd10614,15'd10294,15'd9974,15'd9654,15'd9334,15'd9014,15'd8694,15'd8374,15'd8054,15'd7734,15'd7414,15'd7094,15'd6774,15'd6454,15'd6134,15'd5814,15'd5494,15'd5174,15'd4854,15'd4534,15'd4214,15'd3894,15'd3574,15'd3254,15'd2934,15'd2614,15'd2294,15'd1974,15'd1654,15'd1334,15'd1014,15'd694,15'd374,15'd54,
15'd25335,15'd25015,15'd24695,15'd24375,15'd24055,15'd23735,15'd23415,15'd23095,15'd22775,15'd22455,15'd22135,15'd21815,15'd21495,15'd21175,15'd20855,15'd20535,15'd20215,15'd19895,15'd19575,15'd19255,15'd18935,15'd18615,15'd18295,15'd17975,15'd17655,15'd17335,15'd17015,15'd16695,15'd16375,15'd16055,15'd15735,15'd15415,15'd15095,15'd14775,15'd14455,15'd14135,15'd13815,15'd13495,15'd13175,15'd12855,15'd12535,15'd12215,15'd11895,15'd11575,15'd11255,15'd10935,15'd10615,15'd10295,15'd9975,15'd9655,15'd9335,15'd9015,15'd8695,15'd8375,15'd8055,15'd7735,15'd7415,15'd7095,15'd6775,15'd6455,15'd6135,15'd5815,15'd5495,15'd5175,15'd4855,15'd4535,15'd4215,15'd3895,15'd3575,15'd3255,15'd2935,15'd2615,15'd2295,15'd1975,15'd1655,15'd1335,15'd1015,15'd695,15'd375,15'd55,
15'd25336,15'd25016,15'd24696,15'd24376,15'd24056,15'd23736,15'd23416,15'd23096,15'd22776,15'd22456,15'd22136,15'd21816,15'd21496,15'd21176,15'd20856,15'd20536,15'd20216,15'd19896,15'd19576,15'd19256,15'd18936,15'd18616,15'd18296,15'd17976,15'd17656,15'd17336,15'd17016,15'd16696,15'd16376,15'd16056,15'd15736,15'd15416,15'd15096,15'd14776,15'd14456,15'd14136,15'd13816,15'd13496,15'd13176,15'd12856,15'd12536,15'd12216,15'd11896,15'd11576,15'd11256,15'd10936,15'd10616,15'd10296,15'd9976,15'd9656,15'd9336,15'd9016,15'd8696,15'd8376,15'd8056,15'd7736,15'd7416,15'd7096,15'd6776,15'd6456,15'd6136,15'd5816,15'd5496,15'd5176,15'd4856,15'd4536,15'd4216,15'd3896,15'd3576,15'd3256,15'd2936,15'd2616,15'd2296,15'd1976,15'd1656,15'd1336,15'd1016,15'd696,15'd376,15'd56,
15'd25337,15'd25017,15'd24697,15'd24377,15'd24057,15'd23737,15'd23417,15'd23097,15'd22777,15'd22457,15'd22137,15'd21817,15'd21497,15'd21177,15'd20857,15'd20537,15'd20217,15'd19897,15'd19577,15'd19257,15'd18937,15'd18617,15'd18297,15'd17977,15'd17657,15'd17337,15'd17017,15'd16697,15'd16377,15'd16057,15'd15737,15'd15417,15'd15097,15'd14777,15'd14457,15'd14137,15'd13817,15'd13497,15'd13177,15'd12857,15'd12537,15'd12217,15'd11897,15'd11577,15'd11257,15'd10937,15'd10617,15'd10297,15'd9977,15'd9657,15'd9337,15'd9017,15'd8697,15'd8377,15'd8057,15'd7737,15'd7417,15'd7097,15'd6777,15'd6457,15'd6137,15'd5817,15'd5497,15'd5177,15'd4857,15'd4537,15'd4217,15'd3897,15'd3577,15'd3257,15'd2937,15'd2617,15'd2297,15'd1977,15'd1657,15'd1337,15'd1017,15'd697,15'd377,15'd57,
15'd25338,15'd25018,15'd24698,15'd24378,15'd24058,15'd23738,15'd23418,15'd23098,15'd22778,15'd22458,15'd22138,15'd21818,15'd21498,15'd21178,15'd20858,15'd20538,15'd20218,15'd19898,15'd19578,15'd19258,15'd18938,15'd18618,15'd18298,15'd17978,15'd17658,15'd17338,15'd17018,15'd16698,15'd16378,15'd16058,15'd15738,15'd15418,15'd15098,15'd14778,15'd14458,15'd14138,15'd13818,15'd13498,15'd13178,15'd12858,15'd12538,15'd12218,15'd11898,15'd11578,15'd11258,15'd10938,15'd10618,15'd10298,15'd9978,15'd9658,15'd9338,15'd9018,15'd8698,15'd8378,15'd8058,15'd7738,15'd7418,15'd7098,15'd6778,15'd6458,15'd6138,15'd5818,15'd5498,15'd5178,15'd4858,15'd4538,15'd4218,15'd3898,15'd3578,15'd3258,15'd2938,15'd2618,15'd2298,15'd1978,15'd1658,15'd1338,15'd1018,15'd698,15'd378,15'd58,
15'd25339,15'd25019,15'd24699,15'd24379,15'd24059,15'd23739,15'd23419,15'd23099,15'd22779,15'd22459,15'd22139,15'd21819,15'd21499,15'd21179,15'd20859,15'd20539,15'd20219,15'd19899,15'd19579,15'd19259,15'd18939,15'd18619,15'd18299,15'd17979,15'd17659,15'd17339,15'd17019,15'd16699,15'd16379,15'd16059,15'd15739,15'd15419,15'd15099,15'd14779,15'd14459,15'd14139,15'd13819,15'd13499,15'd13179,15'd12859,15'd12539,15'd12219,15'd11899,15'd11579,15'd11259,15'd10939,15'd10619,15'd10299,15'd9979,15'd9659,15'd9339,15'd9019,15'd8699,15'd8379,15'd8059,15'd7739,15'd7419,15'd7099,15'd6779,15'd6459,15'd6139,15'd5819,15'd5499,15'd5179,15'd4859,15'd4539,15'd4219,15'd3899,15'd3579,15'd3259,15'd2939,15'd2619,15'd2299,15'd1979,15'd1659,15'd1339,15'd1019,15'd699,15'd379,15'd59,
15'd25340,15'd25020,15'd24700,15'd24380,15'd24060,15'd23740,15'd23420,15'd23100,15'd22780,15'd22460,15'd22140,15'd21820,15'd21500,15'd21180,15'd20860,15'd20540,15'd20220,15'd19900,15'd19580,15'd19260,15'd18940,15'd18620,15'd18300,15'd17980,15'd17660,15'd17340,15'd17020,15'd16700,15'd16380,15'd16060,15'd15740,15'd15420,15'd15100,15'd14780,15'd14460,15'd14140,15'd13820,15'd13500,15'd13180,15'd12860,15'd12540,15'd12220,15'd11900,15'd11580,15'd11260,15'd10940,15'd10620,15'd10300,15'd9980,15'd9660,15'd9340,15'd9020,15'd8700,15'd8380,15'd8060,15'd7740,15'd7420,15'd7100,15'd6780,15'd6460,15'd6140,15'd5820,15'd5500,15'd5180,15'd4860,15'd4540,15'd4220,15'd3900,15'd3580,15'd3260,15'd2940,15'd2620,15'd2300,15'd1980,15'd1660,15'd1340,15'd1020,15'd700,15'd380,15'd60,
15'd25341,15'd25021,15'd24701,15'd24381,15'd24061,15'd23741,15'd23421,15'd23101,15'd22781,15'd22461,15'd22141,15'd21821,15'd21501,15'd21181,15'd20861,15'd20541,15'd20221,15'd19901,15'd19581,15'd19261,15'd18941,15'd18621,15'd18301,15'd17981,15'd17661,15'd17341,15'd17021,15'd16701,15'd16381,15'd16061,15'd15741,15'd15421,15'd15101,15'd14781,15'd14461,15'd14141,15'd13821,15'd13501,15'd13181,15'd12861,15'd12541,15'd12221,15'd11901,15'd11581,15'd11261,15'd10941,15'd10621,15'd10301,15'd9981,15'd9661,15'd9341,15'd9021,15'd8701,15'd8381,15'd8061,15'd7741,15'd7421,15'd7101,15'd6781,15'd6461,15'd6141,15'd5821,15'd5501,15'd5181,15'd4861,15'd4541,15'd4221,15'd3901,15'd3581,15'd3261,15'd2941,15'd2621,15'd2301,15'd1981,15'd1661,15'd1341,15'd1021,15'd701,15'd381,15'd61,
15'd25342,15'd25022,15'd24702,15'd24382,15'd24062,15'd23742,15'd23422,15'd23102,15'd22782,15'd22462,15'd22142,15'd21822,15'd21502,15'd21182,15'd20862,15'd20542,15'd20222,15'd19902,15'd19582,15'd19262,15'd18942,15'd18622,15'd18302,15'd17982,15'd17662,15'd17342,15'd17022,15'd16702,15'd16382,15'd16062,15'd15742,15'd15422,15'd15102,15'd14782,15'd14462,15'd14142,15'd13822,15'd13502,15'd13182,15'd12862,15'd12542,15'd12222,15'd11902,15'd11582,15'd11262,15'd10942,15'd10622,15'd10302,15'd9982,15'd9662,15'd9342,15'd9022,15'd8702,15'd8382,15'd8062,15'd7742,15'd7422,15'd7102,15'd6782,15'd6462,15'd6142,15'd5822,15'd5502,15'd5182,15'd4862,15'd4542,15'd4222,15'd3902,15'd3582,15'd3262,15'd2942,15'd2622,15'd2302,15'd1982,15'd1662,15'd1342,15'd1022,15'd702,15'd382,15'd62,
15'd25343,15'd25023,15'd24703,15'd24383,15'd24063,15'd23743,15'd23423,15'd23103,15'd22783,15'd22463,15'd22143,15'd21823,15'd21503,15'd21183,15'd20863,15'd20543,15'd20223,15'd19903,15'd19583,15'd19263,15'd18943,15'd18623,15'd18303,15'd17983,15'd17663,15'd17343,15'd17023,15'd16703,15'd16383,15'd16063,15'd15743,15'd15423,15'd15103,15'd14783,15'd14463,15'd14143,15'd13823,15'd13503,15'd13183,15'd12863,15'd12543,15'd12223,15'd11903,15'd11583,15'd11263,15'd10943,15'd10623,15'd10303,15'd9983,15'd9663,15'd9343,15'd9023,15'd8703,15'd8383,15'd8063,15'd7743,15'd7423,15'd7103,15'd6783,15'd6463,15'd6143,15'd5823,15'd5503,15'd5183,15'd4863,15'd4543,15'd4223,15'd3903,15'd3583,15'd3263,15'd2943,15'd2623,15'd2303,15'd1983,15'd1663,15'd1343,15'd1023,15'd703,15'd383,15'd63,
15'd25344,15'd25024,15'd24704,15'd24384,15'd24064,15'd23744,15'd23424,15'd23104,15'd22784,15'd22464,15'd22144,15'd21824,15'd21504,15'd21184,15'd20864,15'd20544,15'd20224,15'd19904,15'd19584,15'd19264,15'd18944,15'd18624,15'd18304,15'd17984,15'd17664,15'd17344,15'd17024,15'd16704,15'd16384,15'd16064,15'd15744,15'd15424,15'd15104,15'd14784,15'd14464,15'd14144,15'd13824,15'd13504,15'd13184,15'd12864,15'd12544,15'd12224,15'd11904,15'd11584,15'd11264,15'd10944,15'd10624,15'd10304,15'd9984,15'd9664,15'd9344,15'd9024,15'd8704,15'd8384,15'd8064,15'd7744,15'd7424,15'd7104,15'd6784,15'd6464,15'd6144,15'd5824,15'd5504,15'd5184,15'd4864,15'd4544,15'd4224,15'd3904,15'd3584,15'd3264,15'd2944,15'd2624,15'd2304,15'd1984,15'd1664,15'd1344,15'd1024,15'd704,15'd384,15'd64,
15'd25345,15'd25025,15'd24705,15'd24385,15'd24065,15'd23745,15'd23425,15'd23105,15'd22785,15'd22465,15'd22145,15'd21825,15'd21505,15'd21185,15'd20865,15'd20545,15'd20225,15'd19905,15'd19585,15'd19265,15'd18945,15'd18625,15'd18305,15'd17985,15'd17665,15'd17345,15'd17025,15'd16705,15'd16385,15'd16065,15'd15745,15'd15425,15'd15105,15'd14785,15'd14465,15'd14145,15'd13825,15'd13505,15'd13185,15'd12865,15'd12545,15'd12225,15'd11905,15'd11585,15'd11265,15'd10945,15'd10625,15'd10305,15'd9985,15'd9665,15'd9345,15'd9025,15'd8705,15'd8385,15'd8065,15'd7745,15'd7425,15'd7105,15'd6785,15'd6465,15'd6145,15'd5825,15'd5505,15'd5185,15'd4865,15'd4545,15'd4225,15'd3905,15'd3585,15'd3265,15'd2945,15'd2625,15'd2305,15'd1985,15'd1665,15'd1345,15'd1025,15'd705,15'd385,15'd65,
15'd25346,15'd25026,15'd24706,15'd24386,15'd24066,15'd23746,15'd23426,15'd23106,15'd22786,15'd22466,15'd22146,15'd21826,15'd21506,15'd21186,15'd20866,15'd20546,15'd20226,15'd19906,15'd19586,15'd19266,15'd18946,15'd18626,15'd18306,15'd17986,15'd17666,15'd17346,15'd17026,15'd16706,15'd16386,15'd16066,15'd15746,15'd15426,15'd15106,15'd14786,15'd14466,15'd14146,15'd13826,15'd13506,15'd13186,15'd12866,15'd12546,15'd12226,15'd11906,15'd11586,15'd11266,15'd10946,15'd10626,15'd10306,15'd9986,15'd9666,15'd9346,15'd9026,15'd8706,15'd8386,15'd8066,15'd7746,15'd7426,15'd7106,15'd6786,15'd6466,15'd6146,15'd5826,15'd5506,15'd5186,15'd4866,15'd4546,15'd4226,15'd3906,15'd3586,15'd3266,15'd2946,15'd2626,15'd2306,15'd1986,15'd1666,15'd1346,15'd1026,15'd706,15'd386,15'd66,
15'd25347,15'd25027,15'd24707,15'd24387,15'd24067,15'd23747,15'd23427,15'd23107,15'd22787,15'd22467,15'd22147,15'd21827,15'd21507,15'd21187,15'd20867,15'd20547,15'd20227,15'd19907,15'd19587,15'd19267,15'd18947,15'd18627,15'd18307,15'd17987,15'd17667,15'd17347,15'd17027,15'd16707,15'd16387,15'd16067,15'd15747,15'd15427,15'd15107,15'd14787,15'd14467,15'd14147,15'd13827,15'd13507,15'd13187,15'd12867,15'd12547,15'd12227,15'd11907,15'd11587,15'd11267,15'd10947,15'd10627,15'd10307,15'd9987,15'd9667,15'd9347,15'd9027,15'd8707,15'd8387,15'd8067,15'd7747,15'd7427,15'd7107,15'd6787,15'd6467,15'd6147,15'd5827,15'd5507,15'd5187,15'd4867,15'd4547,15'd4227,15'd3907,15'd3587,15'd3267,15'd2947,15'd2627,15'd2307,15'd1987,15'd1667,15'd1347,15'd1027,15'd707,15'd387,15'd67,
15'd25348,15'd25028,15'd24708,15'd24388,15'd24068,15'd23748,15'd23428,15'd23108,15'd22788,15'd22468,15'd22148,15'd21828,15'd21508,15'd21188,15'd20868,15'd20548,15'd20228,15'd19908,15'd19588,15'd19268,15'd18948,15'd18628,15'd18308,15'd17988,15'd17668,15'd17348,15'd17028,15'd16708,15'd16388,15'd16068,15'd15748,15'd15428,15'd15108,15'd14788,15'd14468,15'd14148,15'd13828,15'd13508,15'd13188,15'd12868,15'd12548,15'd12228,15'd11908,15'd11588,15'd11268,15'd10948,15'd10628,15'd10308,15'd9988,15'd9668,15'd9348,15'd9028,15'd8708,15'd8388,15'd8068,15'd7748,15'd7428,15'd7108,15'd6788,15'd6468,15'd6148,15'd5828,15'd5508,15'd5188,15'd4868,15'd4548,15'd4228,15'd3908,15'd3588,15'd3268,15'd2948,15'd2628,15'd2308,15'd1988,15'd1668,15'd1348,15'd1028,15'd708,15'd388,15'd68,
15'd25349,15'd25029,15'd24709,15'd24389,15'd24069,15'd23749,15'd23429,15'd23109,15'd22789,15'd22469,15'd22149,15'd21829,15'd21509,15'd21189,15'd20869,15'd20549,15'd20229,15'd19909,15'd19589,15'd19269,15'd18949,15'd18629,15'd18309,15'd17989,15'd17669,15'd17349,15'd17029,15'd16709,15'd16389,15'd16069,15'd15749,15'd15429,15'd15109,15'd14789,15'd14469,15'd14149,15'd13829,15'd13509,15'd13189,15'd12869,15'd12549,15'd12229,15'd11909,15'd11589,15'd11269,15'd10949,15'd10629,15'd10309,15'd9989,15'd9669,15'd9349,15'd9029,15'd8709,15'd8389,15'd8069,15'd7749,15'd7429,15'd7109,15'd6789,15'd6469,15'd6149,15'd5829,15'd5509,15'd5189,15'd4869,15'd4549,15'd4229,15'd3909,15'd3589,15'd3269,15'd2949,15'd2629,15'd2309,15'd1989,15'd1669,15'd1349,15'd1029,15'd709,15'd389,15'd69,
15'd25350,15'd25030,15'd24710,15'd24390,15'd24070,15'd23750,15'd23430,15'd23110,15'd22790,15'd22470,15'd22150,15'd21830,15'd21510,15'd21190,15'd20870,15'd20550,15'd20230,15'd19910,15'd19590,15'd19270,15'd18950,15'd18630,15'd18310,15'd17990,15'd17670,15'd17350,15'd17030,15'd16710,15'd16390,15'd16070,15'd15750,15'd15430,15'd15110,15'd14790,15'd14470,15'd14150,15'd13830,15'd13510,15'd13190,15'd12870,15'd12550,15'd12230,15'd11910,15'd11590,15'd11270,15'd10950,15'd10630,15'd10310,15'd9990,15'd9670,15'd9350,15'd9030,15'd8710,15'd8390,15'd8070,15'd7750,15'd7430,15'd7110,15'd6790,15'd6470,15'd6150,15'd5830,15'd5510,15'd5190,15'd4870,15'd4550,15'd4230,15'd3910,15'd3590,15'd3270,15'd2950,15'd2630,15'd2310,15'd1990,15'd1670,15'd1350,15'd1030,15'd710,15'd390,15'd70,
15'd25351,15'd25031,15'd24711,15'd24391,15'd24071,15'd23751,15'd23431,15'd23111,15'd22791,15'd22471,15'd22151,15'd21831,15'd21511,15'd21191,15'd20871,15'd20551,15'd20231,15'd19911,15'd19591,15'd19271,15'd18951,15'd18631,15'd18311,15'd17991,15'd17671,15'd17351,15'd17031,15'd16711,15'd16391,15'd16071,15'd15751,15'd15431,15'd15111,15'd14791,15'd14471,15'd14151,15'd13831,15'd13511,15'd13191,15'd12871,15'd12551,15'd12231,15'd11911,15'd11591,15'd11271,15'd10951,15'd10631,15'd10311,15'd9991,15'd9671,15'd9351,15'd9031,15'd8711,15'd8391,15'd8071,15'd7751,15'd7431,15'd7111,15'd6791,15'd6471,15'd6151,15'd5831,15'd5511,15'd5191,15'd4871,15'd4551,15'd4231,15'd3911,15'd3591,15'd3271,15'd2951,15'd2631,15'd2311,15'd1991,15'd1671,15'd1351,15'd1031,15'd711,15'd391,15'd71,
15'd25352,15'd25032,15'd24712,15'd24392,15'd24072,15'd23752,15'd23432,15'd23112,15'd22792,15'd22472,15'd22152,15'd21832,15'd21512,15'd21192,15'd20872,15'd20552,15'd20232,15'd19912,15'd19592,15'd19272,15'd18952,15'd18632,15'd18312,15'd17992,15'd17672,15'd17352,15'd17032,15'd16712,15'd16392,15'd16072,15'd15752,15'd15432,15'd15112,15'd14792,15'd14472,15'd14152,15'd13832,15'd13512,15'd13192,15'd12872,15'd12552,15'd12232,15'd11912,15'd11592,15'd11272,15'd10952,15'd10632,15'd10312,15'd9992,15'd9672,15'd9352,15'd9032,15'd8712,15'd8392,15'd8072,15'd7752,15'd7432,15'd7112,15'd6792,15'd6472,15'd6152,15'd5832,15'd5512,15'd5192,15'd4872,15'd4552,15'd4232,15'd3912,15'd3592,15'd3272,15'd2952,15'd2632,15'd2312,15'd1992,15'd1672,15'd1352,15'd1032,15'd712,15'd392,15'd72,
15'd25353,15'd25033,15'd24713,15'd24393,15'd24073,15'd23753,15'd23433,15'd23113,15'd22793,15'd22473,15'd22153,15'd21833,15'd21513,15'd21193,15'd20873,15'd20553,15'd20233,15'd19913,15'd19593,15'd19273,15'd18953,15'd18633,15'd18313,15'd17993,15'd17673,15'd17353,15'd17033,15'd16713,15'd16393,15'd16073,15'd15753,15'd15433,15'd15113,15'd14793,15'd14473,15'd14153,15'd13833,15'd13513,15'd13193,15'd12873,15'd12553,15'd12233,15'd11913,15'd11593,15'd11273,15'd10953,15'd10633,15'd10313,15'd9993,15'd9673,15'd9353,15'd9033,15'd8713,15'd8393,15'd8073,15'd7753,15'd7433,15'd7113,15'd6793,15'd6473,15'd6153,15'd5833,15'd5513,15'd5193,15'd4873,15'd4553,15'd4233,15'd3913,15'd3593,15'd3273,15'd2953,15'd2633,15'd2313,15'd1993,15'd1673,15'd1353,15'd1033,15'd713,15'd393,15'd73,
15'd25354,15'd25034,15'd24714,15'd24394,15'd24074,15'd23754,15'd23434,15'd23114,15'd22794,15'd22474,15'd22154,15'd21834,15'd21514,15'd21194,15'd20874,15'd20554,15'd20234,15'd19914,15'd19594,15'd19274,15'd18954,15'd18634,15'd18314,15'd17994,15'd17674,15'd17354,15'd17034,15'd16714,15'd16394,15'd16074,15'd15754,15'd15434,15'd15114,15'd14794,15'd14474,15'd14154,15'd13834,15'd13514,15'd13194,15'd12874,15'd12554,15'd12234,15'd11914,15'd11594,15'd11274,15'd10954,15'd10634,15'd10314,15'd9994,15'd9674,15'd9354,15'd9034,15'd8714,15'd8394,15'd8074,15'd7754,15'd7434,15'd7114,15'd6794,15'd6474,15'd6154,15'd5834,15'd5514,15'd5194,15'd4874,15'd4554,15'd4234,15'd3914,15'd3594,15'd3274,15'd2954,15'd2634,15'd2314,15'd1994,15'd1674,15'd1354,15'd1034,15'd714,15'd394,15'd74,
15'd25355,15'd25035,15'd24715,15'd24395,15'd24075,15'd23755,15'd23435,15'd23115,15'd22795,15'd22475,15'd22155,15'd21835,15'd21515,15'd21195,15'd20875,15'd20555,15'd20235,15'd19915,15'd19595,15'd19275,15'd18955,15'd18635,15'd18315,15'd17995,15'd17675,15'd17355,15'd17035,15'd16715,15'd16395,15'd16075,15'd15755,15'd15435,15'd15115,15'd14795,15'd14475,15'd14155,15'd13835,15'd13515,15'd13195,15'd12875,15'd12555,15'd12235,15'd11915,15'd11595,15'd11275,15'd10955,15'd10635,15'd10315,15'd9995,15'd9675,15'd9355,15'd9035,15'd8715,15'd8395,15'd8075,15'd7755,15'd7435,15'd7115,15'd6795,15'd6475,15'd6155,15'd5835,15'd5515,15'd5195,15'd4875,15'd4555,15'd4235,15'd3915,15'd3595,15'd3275,15'd2955,15'd2635,15'd2315,15'd1995,15'd1675,15'd1355,15'd1035,15'd715,15'd395,15'd75,
15'd25356,15'd25036,15'd24716,15'd24396,15'd24076,15'd23756,15'd23436,15'd23116,15'd22796,15'd22476,15'd22156,15'd21836,15'd21516,15'd21196,15'd20876,15'd20556,15'd20236,15'd19916,15'd19596,15'd19276,15'd18956,15'd18636,15'd18316,15'd17996,15'd17676,15'd17356,15'd17036,15'd16716,15'd16396,15'd16076,15'd15756,15'd15436,15'd15116,15'd14796,15'd14476,15'd14156,15'd13836,15'd13516,15'd13196,15'd12876,15'd12556,15'd12236,15'd11916,15'd11596,15'd11276,15'd10956,15'd10636,15'd10316,15'd9996,15'd9676,15'd9356,15'd9036,15'd8716,15'd8396,15'd8076,15'd7756,15'd7436,15'd7116,15'd6796,15'd6476,15'd6156,15'd5836,15'd5516,15'd5196,15'd4876,15'd4556,15'd4236,15'd3916,15'd3596,15'd3276,15'd2956,15'd2636,15'd2316,15'd1996,15'd1676,15'd1356,15'd1036,15'd716,15'd396,15'd76,
15'd25357,15'd25037,15'd24717,15'd24397,15'd24077,15'd23757,15'd23437,15'd23117,15'd22797,15'd22477,15'd22157,15'd21837,15'd21517,15'd21197,15'd20877,15'd20557,15'd20237,15'd19917,15'd19597,15'd19277,15'd18957,15'd18637,15'd18317,15'd17997,15'd17677,15'd17357,15'd17037,15'd16717,15'd16397,15'd16077,15'd15757,15'd15437,15'd15117,15'd14797,15'd14477,15'd14157,15'd13837,15'd13517,15'd13197,15'd12877,15'd12557,15'd12237,15'd11917,15'd11597,15'd11277,15'd10957,15'd10637,15'd10317,15'd9997,15'd9677,15'd9357,15'd9037,15'd8717,15'd8397,15'd8077,15'd7757,15'd7437,15'd7117,15'd6797,15'd6477,15'd6157,15'd5837,15'd5517,15'd5197,15'd4877,15'd4557,15'd4237,15'd3917,15'd3597,15'd3277,15'd2957,15'd2637,15'd2317,15'd1997,15'd1677,15'd1357,15'd1037,15'd717,15'd397,15'd77,
15'd25358,15'd25038,15'd24718,15'd24398,15'd24078,15'd23758,15'd23438,15'd23118,15'd22798,15'd22478,15'd22158,15'd21838,15'd21518,15'd21198,15'd20878,15'd20558,15'd20238,15'd19918,15'd19598,15'd19278,15'd18958,15'd18638,15'd18318,15'd17998,15'd17678,15'd17358,15'd17038,15'd16718,15'd16398,15'd16078,15'd15758,15'd15438,15'd15118,15'd14798,15'd14478,15'd14158,15'd13838,15'd13518,15'd13198,15'd12878,15'd12558,15'd12238,15'd11918,15'd11598,15'd11278,15'd10958,15'd10638,15'd10318,15'd9998,15'd9678,15'd9358,15'd9038,15'd8718,15'd8398,15'd8078,15'd7758,15'd7438,15'd7118,15'd6798,15'd6478,15'd6158,15'd5838,15'd5518,15'd5198,15'd4878,15'd4558,15'd4238,15'd3918,15'd3598,15'd3278,15'd2958,15'd2638,15'd2318,15'd1998,15'd1678,15'd1358,15'd1038,15'd718,15'd398,15'd78,
15'd25359,15'd25039,15'd24719,15'd24399,15'd24079,15'd23759,15'd23439,15'd23119,15'd22799,15'd22479,15'd22159,15'd21839,15'd21519,15'd21199,15'd20879,15'd20559,15'd20239,15'd19919,15'd19599,15'd19279,15'd18959,15'd18639,15'd18319,15'd17999,15'd17679,15'd17359,15'd17039,15'd16719,15'd16399,15'd16079,15'd15759,15'd15439,15'd15119,15'd14799,15'd14479,15'd14159,15'd13839,15'd13519,15'd13199,15'd12879,15'd12559,15'd12239,15'd11919,15'd11599,15'd11279,15'd10959,15'd10639,15'd10319,15'd9999,15'd9679,15'd9359,15'd9039,15'd8719,15'd8399,15'd8079,15'd7759,15'd7439,15'd7119,15'd6799,15'd6479,15'd6159,15'd5839,15'd5519,15'd5199,15'd4879,15'd4559,15'd4239,15'd3919,15'd3599,15'd3279,15'd2959,15'd2639,15'd2319,15'd1999,15'd1679,15'd1359,15'd1039,15'd719,15'd399,15'd79};
parameter [14:0] state_2 [0:6399] = {
15'd25359,15'd25358,15'd25357,15'd25356,15'd25355,15'd25354,15'd25353,15'd25352,15'd25351,15'd25350,15'd25349,15'd25348,15'd25347,15'd25346,15'd25345,15'd25344,15'd25343,15'd25342,15'd25341,15'd25340,15'd25339,15'd25338,15'd25337,15'd25336,15'd25335,15'd25334,15'd25333,15'd25332,15'd25331,15'd25330,15'd25329,15'd25328,15'd25327,15'd25326,15'd25325,15'd25324,15'd25323,15'd25322,15'd25321,15'd25320,15'd25319,15'd25318,15'd25317,15'd25316,15'd25315,15'd25314,15'd25313,15'd25312,15'd25311,15'd25310,15'd25309,15'd25308,15'd25307,15'd25306,15'd25305,15'd25304,15'd25303,15'd25302,15'd25301,15'd25300,15'd25299,15'd25298,15'd25297,15'd25296,15'd25295,15'd25294,15'd25293,15'd25292,15'd25291,15'd25290,15'd25289,15'd25288,15'd25287,15'd25286,15'd25285,15'd25284,15'd25283,15'd25282,15'd25281,15'd25280,
15'd25039,15'd25038,15'd25037,15'd25036,15'd25035,15'd25034,15'd25033,15'd25032,15'd25031,15'd25030,15'd25029,15'd25028,15'd25027,15'd25026,15'd25025,15'd25024,15'd25023,15'd25022,15'd25021,15'd25020,15'd25019,15'd25018,15'd25017,15'd25016,15'd25015,15'd25014,15'd25013,15'd25012,15'd25011,15'd25010,15'd25009,15'd25008,15'd25007,15'd25006,15'd25005,15'd25004,15'd25003,15'd25002,15'd25001,15'd25000,15'd24999,15'd24998,15'd24997,15'd24996,15'd24995,15'd24994,15'd24993,15'd24992,15'd24991,15'd24990,15'd24989,15'd24988,15'd24987,15'd24986,15'd24985,15'd24984,15'd24983,15'd24982,15'd24981,15'd24980,15'd24979,15'd24978,15'd24977,15'd24976,15'd24975,15'd24974,15'd24973,15'd24972,15'd24971,15'd24970,15'd24969,15'd24968,15'd24967,15'd24966,15'd24965,15'd24964,15'd24963,15'd24962,15'd24961,15'd24960,
15'd24719,15'd24718,15'd24717,15'd24716,15'd24715,15'd24714,15'd24713,15'd24712,15'd24711,15'd24710,15'd24709,15'd24708,15'd24707,15'd24706,15'd24705,15'd24704,15'd24703,15'd24702,15'd24701,15'd24700,15'd24699,15'd24698,15'd24697,15'd24696,15'd24695,15'd24694,15'd24693,15'd24692,15'd24691,15'd24690,15'd24689,15'd24688,15'd24687,15'd24686,15'd24685,15'd24684,15'd24683,15'd24682,15'd24681,15'd24680,15'd24679,15'd24678,15'd24677,15'd24676,15'd24675,15'd24674,15'd24673,15'd24672,15'd24671,15'd24670,15'd24669,15'd24668,15'd24667,15'd24666,15'd24665,15'd24664,15'd24663,15'd24662,15'd24661,15'd24660,15'd24659,15'd24658,15'd24657,15'd24656,15'd24655,15'd24654,15'd24653,15'd24652,15'd24651,15'd24650,15'd24649,15'd24648,15'd24647,15'd24646,15'd24645,15'd24644,15'd24643,15'd24642,15'd24641,15'd24640,
15'd24399,15'd24398,15'd24397,15'd24396,15'd24395,15'd24394,15'd24393,15'd24392,15'd24391,15'd24390,15'd24389,15'd24388,15'd24387,15'd24386,15'd24385,15'd24384,15'd24383,15'd24382,15'd24381,15'd24380,15'd24379,15'd24378,15'd24377,15'd24376,15'd24375,15'd24374,15'd24373,15'd24372,15'd24371,15'd24370,15'd24369,15'd24368,15'd24367,15'd24366,15'd24365,15'd24364,15'd24363,15'd24362,15'd24361,15'd24360,15'd24359,15'd24358,15'd24357,15'd24356,15'd24355,15'd24354,15'd24353,15'd24352,15'd24351,15'd24350,15'd24349,15'd24348,15'd24347,15'd24346,15'd24345,15'd24344,15'd24343,15'd24342,15'd24341,15'd24340,15'd24339,15'd24338,15'd24337,15'd24336,15'd24335,15'd24334,15'd24333,15'd24332,15'd24331,15'd24330,15'd24329,15'd24328,15'd24327,15'd24326,15'd24325,15'd24324,15'd24323,15'd24322,15'd24321,15'd24320,
15'd24079,15'd24078,15'd24077,15'd24076,15'd24075,15'd24074,15'd24073,15'd24072,15'd24071,15'd24070,15'd24069,15'd24068,15'd24067,15'd24066,15'd24065,15'd24064,15'd24063,15'd24062,15'd24061,15'd24060,15'd24059,15'd24058,15'd24057,15'd24056,15'd24055,15'd24054,15'd24053,15'd24052,15'd24051,15'd24050,15'd24049,15'd24048,15'd24047,15'd24046,15'd24045,15'd24044,15'd24043,15'd24042,15'd24041,15'd24040,15'd24039,15'd24038,15'd24037,15'd24036,15'd24035,15'd24034,15'd24033,15'd24032,15'd24031,15'd24030,15'd24029,15'd24028,15'd24027,15'd24026,15'd24025,15'd24024,15'd24023,15'd24022,15'd24021,15'd24020,15'd24019,15'd24018,15'd24017,15'd24016,15'd24015,15'd24014,15'd24013,15'd24012,15'd24011,15'd24010,15'd24009,15'd24008,15'd24007,15'd24006,15'd24005,15'd24004,15'd24003,15'd24002,15'd24001,15'd24000,
15'd23759,15'd23758,15'd23757,15'd23756,15'd23755,15'd23754,15'd23753,15'd23752,15'd23751,15'd23750,15'd23749,15'd23748,15'd23747,15'd23746,15'd23745,15'd23744,15'd23743,15'd23742,15'd23741,15'd23740,15'd23739,15'd23738,15'd23737,15'd23736,15'd23735,15'd23734,15'd23733,15'd23732,15'd23731,15'd23730,15'd23729,15'd23728,15'd23727,15'd23726,15'd23725,15'd23724,15'd23723,15'd23722,15'd23721,15'd23720,15'd23719,15'd23718,15'd23717,15'd23716,15'd23715,15'd23714,15'd23713,15'd23712,15'd23711,15'd23710,15'd23709,15'd23708,15'd23707,15'd23706,15'd23705,15'd23704,15'd23703,15'd23702,15'd23701,15'd23700,15'd23699,15'd23698,15'd23697,15'd23696,15'd23695,15'd23694,15'd23693,15'd23692,15'd23691,15'd23690,15'd23689,15'd23688,15'd23687,15'd23686,15'd23685,15'd23684,15'd23683,15'd23682,15'd23681,15'd23680,
15'd23439,15'd23438,15'd23437,15'd23436,15'd23435,15'd23434,15'd23433,15'd23432,15'd23431,15'd23430,15'd23429,15'd23428,15'd23427,15'd23426,15'd23425,15'd23424,15'd23423,15'd23422,15'd23421,15'd23420,15'd23419,15'd23418,15'd23417,15'd23416,15'd23415,15'd23414,15'd23413,15'd23412,15'd23411,15'd23410,15'd23409,15'd23408,15'd23407,15'd23406,15'd23405,15'd23404,15'd23403,15'd23402,15'd23401,15'd23400,15'd23399,15'd23398,15'd23397,15'd23396,15'd23395,15'd23394,15'd23393,15'd23392,15'd23391,15'd23390,15'd23389,15'd23388,15'd23387,15'd23386,15'd23385,15'd23384,15'd23383,15'd23382,15'd23381,15'd23380,15'd23379,15'd23378,15'd23377,15'd23376,15'd23375,15'd23374,15'd23373,15'd23372,15'd23371,15'd23370,15'd23369,15'd23368,15'd23367,15'd23366,15'd23365,15'd23364,15'd23363,15'd23362,15'd23361,15'd23360,
15'd23119,15'd23118,15'd23117,15'd23116,15'd23115,15'd23114,15'd23113,15'd23112,15'd23111,15'd23110,15'd23109,15'd23108,15'd23107,15'd23106,15'd23105,15'd23104,15'd23103,15'd23102,15'd23101,15'd23100,15'd23099,15'd23098,15'd23097,15'd23096,15'd23095,15'd23094,15'd23093,15'd23092,15'd23091,15'd23090,15'd23089,15'd23088,15'd23087,15'd23086,15'd23085,15'd23084,15'd23083,15'd23082,15'd23081,15'd23080,15'd23079,15'd23078,15'd23077,15'd23076,15'd23075,15'd23074,15'd23073,15'd23072,15'd23071,15'd23070,15'd23069,15'd23068,15'd23067,15'd23066,15'd23065,15'd23064,15'd23063,15'd23062,15'd23061,15'd23060,15'd23059,15'd23058,15'd23057,15'd23056,15'd23055,15'd23054,15'd23053,15'd23052,15'd23051,15'd23050,15'd23049,15'd23048,15'd23047,15'd23046,15'd23045,15'd23044,15'd23043,15'd23042,15'd23041,15'd23040,
15'd22799,15'd22798,15'd22797,15'd22796,15'd22795,15'd22794,15'd22793,15'd22792,15'd22791,15'd22790,15'd22789,15'd22788,15'd22787,15'd22786,15'd22785,15'd22784,15'd22783,15'd22782,15'd22781,15'd22780,15'd22779,15'd22778,15'd22777,15'd22776,15'd22775,15'd22774,15'd22773,15'd22772,15'd22771,15'd22770,15'd22769,15'd22768,15'd22767,15'd22766,15'd22765,15'd22764,15'd22763,15'd22762,15'd22761,15'd22760,15'd22759,15'd22758,15'd22757,15'd22756,15'd22755,15'd22754,15'd22753,15'd22752,15'd22751,15'd22750,15'd22749,15'd22748,15'd22747,15'd22746,15'd22745,15'd22744,15'd22743,15'd22742,15'd22741,15'd22740,15'd22739,15'd22738,15'd22737,15'd22736,15'd22735,15'd22734,15'd22733,15'd22732,15'd22731,15'd22730,15'd22729,15'd22728,15'd22727,15'd22726,15'd22725,15'd22724,15'd22723,15'd22722,15'd22721,15'd22720,
15'd22479,15'd22478,15'd22477,15'd22476,15'd22475,15'd22474,15'd22473,15'd22472,15'd22471,15'd22470,15'd22469,15'd22468,15'd22467,15'd22466,15'd22465,15'd22464,15'd22463,15'd22462,15'd22461,15'd22460,15'd22459,15'd22458,15'd22457,15'd22456,15'd22455,15'd22454,15'd22453,15'd22452,15'd22451,15'd22450,15'd22449,15'd22448,15'd22447,15'd22446,15'd22445,15'd22444,15'd22443,15'd22442,15'd22441,15'd22440,15'd22439,15'd22438,15'd22437,15'd22436,15'd22435,15'd22434,15'd22433,15'd22432,15'd22431,15'd22430,15'd22429,15'd22428,15'd22427,15'd22426,15'd22425,15'd22424,15'd22423,15'd22422,15'd22421,15'd22420,15'd22419,15'd22418,15'd22417,15'd22416,15'd22415,15'd22414,15'd22413,15'd22412,15'd22411,15'd22410,15'd22409,15'd22408,15'd22407,15'd22406,15'd22405,15'd22404,15'd22403,15'd22402,15'd22401,15'd22400,
15'd22159,15'd22158,15'd22157,15'd22156,15'd22155,15'd22154,15'd22153,15'd22152,15'd22151,15'd22150,15'd22149,15'd22148,15'd22147,15'd22146,15'd22145,15'd22144,15'd22143,15'd22142,15'd22141,15'd22140,15'd22139,15'd22138,15'd22137,15'd22136,15'd22135,15'd22134,15'd22133,15'd22132,15'd22131,15'd22130,15'd22129,15'd22128,15'd22127,15'd22126,15'd22125,15'd22124,15'd22123,15'd22122,15'd22121,15'd22120,15'd22119,15'd22118,15'd22117,15'd22116,15'd22115,15'd22114,15'd22113,15'd22112,15'd22111,15'd22110,15'd22109,15'd22108,15'd22107,15'd22106,15'd22105,15'd22104,15'd22103,15'd22102,15'd22101,15'd22100,15'd22099,15'd22098,15'd22097,15'd22096,15'd22095,15'd22094,15'd22093,15'd22092,15'd22091,15'd22090,15'd22089,15'd22088,15'd22087,15'd22086,15'd22085,15'd22084,15'd22083,15'd22082,15'd22081,15'd22080,
15'd21839,15'd21838,15'd21837,15'd21836,15'd21835,15'd21834,15'd21833,15'd21832,15'd21831,15'd21830,15'd21829,15'd21828,15'd21827,15'd21826,15'd21825,15'd21824,15'd21823,15'd21822,15'd21821,15'd21820,15'd21819,15'd21818,15'd21817,15'd21816,15'd21815,15'd21814,15'd21813,15'd21812,15'd21811,15'd21810,15'd21809,15'd21808,15'd21807,15'd21806,15'd21805,15'd21804,15'd21803,15'd21802,15'd21801,15'd21800,15'd21799,15'd21798,15'd21797,15'd21796,15'd21795,15'd21794,15'd21793,15'd21792,15'd21791,15'd21790,15'd21789,15'd21788,15'd21787,15'd21786,15'd21785,15'd21784,15'd21783,15'd21782,15'd21781,15'd21780,15'd21779,15'd21778,15'd21777,15'd21776,15'd21775,15'd21774,15'd21773,15'd21772,15'd21771,15'd21770,15'd21769,15'd21768,15'd21767,15'd21766,15'd21765,15'd21764,15'd21763,15'd21762,15'd21761,15'd21760,
15'd21519,15'd21518,15'd21517,15'd21516,15'd21515,15'd21514,15'd21513,15'd21512,15'd21511,15'd21510,15'd21509,15'd21508,15'd21507,15'd21506,15'd21505,15'd21504,15'd21503,15'd21502,15'd21501,15'd21500,15'd21499,15'd21498,15'd21497,15'd21496,15'd21495,15'd21494,15'd21493,15'd21492,15'd21491,15'd21490,15'd21489,15'd21488,15'd21487,15'd21486,15'd21485,15'd21484,15'd21483,15'd21482,15'd21481,15'd21480,15'd21479,15'd21478,15'd21477,15'd21476,15'd21475,15'd21474,15'd21473,15'd21472,15'd21471,15'd21470,15'd21469,15'd21468,15'd21467,15'd21466,15'd21465,15'd21464,15'd21463,15'd21462,15'd21461,15'd21460,15'd21459,15'd21458,15'd21457,15'd21456,15'd21455,15'd21454,15'd21453,15'd21452,15'd21451,15'd21450,15'd21449,15'd21448,15'd21447,15'd21446,15'd21445,15'd21444,15'd21443,15'd21442,15'd21441,15'd21440,
15'd21199,15'd21198,15'd21197,15'd21196,15'd21195,15'd21194,15'd21193,15'd21192,15'd21191,15'd21190,15'd21189,15'd21188,15'd21187,15'd21186,15'd21185,15'd21184,15'd21183,15'd21182,15'd21181,15'd21180,15'd21179,15'd21178,15'd21177,15'd21176,15'd21175,15'd21174,15'd21173,15'd21172,15'd21171,15'd21170,15'd21169,15'd21168,15'd21167,15'd21166,15'd21165,15'd21164,15'd21163,15'd21162,15'd21161,15'd21160,15'd21159,15'd21158,15'd21157,15'd21156,15'd21155,15'd21154,15'd21153,15'd21152,15'd21151,15'd21150,15'd21149,15'd21148,15'd21147,15'd21146,15'd21145,15'd21144,15'd21143,15'd21142,15'd21141,15'd21140,15'd21139,15'd21138,15'd21137,15'd21136,15'd21135,15'd21134,15'd21133,15'd21132,15'd21131,15'd21130,15'd21129,15'd21128,15'd21127,15'd21126,15'd21125,15'd21124,15'd21123,15'd21122,15'd21121,15'd21120,
15'd20879,15'd20878,15'd20877,15'd20876,15'd20875,15'd20874,15'd20873,15'd20872,15'd20871,15'd20870,15'd20869,15'd20868,15'd20867,15'd20866,15'd20865,15'd20864,15'd20863,15'd20862,15'd20861,15'd20860,15'd20859,15'd20858,15'd20857,15'd20856,15'd20855,15'd20854,15'd20853,15'd20852,15'd20851,15'd20850,15'd20849,15'd20848,15'd20847,15'd20846,15'd20845,15'd20844,15'd20843,15'd20842,15'd20841,15'd20840,15'd20839,15'd20838,15'd20837,15'd20836,15'd20835,15'd20834,15'd20833,15'd20832,15'd20831,15'd20830,15'd20829,15'd20828,15'd20827,15'd20826,15'd20825,15'd20824,15'd20823,15'd20822,15'd20821,15'd20820,15'd20819,15'd20818,15'd20817,15'd20816,15'd20815,15'd20814,15'd20813,15'd20812,15'd20811,15'd20810,15'd20809,15'd20808,15'd20807,15'd20806,15'd20805,15'd20804,15'd20803,15'd20802,15'd20801,15'd20800,
15'd20559,15'd20558,15'd20557,15'd20556,15'd20555,15'd20554,15'd20553,15'd20552,15'd20551,15'd20550,15'd20549,15'd20548,15'd20547,15'd20546,15'd20545,15'd20544,15'd20543,15'd20542,15'd20541,15'd20540,15'd20539,15'd20538,15'd20537,15'd20536,15'd20535,15'd20534,15'd20533,15'd20532,15'd20531,15'd20530,15'd20529,15'd20528,15'd20527,15'd20526,15'd20525,15'd20524,15'd20523,15'd20522,15'd20521,15'd20520,15'd20519,15'd20518,15'd20517,15'd20516,15'd20515,15'd20514,15'd20513,15'd20512,15'd20511,15'd20510,15'd20509,15'd20508,15'd20507,15'd20506,15'd20505,15'd20504,15'd20503,15'd20502,15'd20501,15'd20500,15'd20499,15'd20498,15'd20497,15'd20496,15'd20495,15'd20494,15'd20493,15'd20492,15'd20491,15'd20490,15'd20489,15'd20488,15'd20487,15'd20486,15'd20485,15'd20484,15'd20483,15'd20482,15'd20481,15'd20480,
15'd20239,15'd20238,15'd20237,15'd20236,15'd20235,15'd20234,15'd20233,15'd20232,15'd20231,15'd20230,15'd20229,15'd20228,15'd20227,15'd20226,15'd20225,15'd20224,15'd20223,15'd20222,15'd20221,15'd20220,15'd20219,15'd20218,15'd20217,15'd20216,15'd20215,15'd20214,15'd20213,15'd20212,15'd20211,15'd20210,15'd20209,15'd20208,15'd20207,15'd20206,15'd20205,15'd20204,15'd20203,15'd20202,15'd20201,15'd20200,15'd20199,15'd20198,15'd20197,15'd20196,15'd20195,15'd20194,15'd20193,15'd20192,15'd20191,15'd20190,15'd20189,15'd20188,15'd20187,15'd20186,15'd20185,15'd20184,15'd20183,15'd20182,15'd20181,15'd20180,15'd20179,15'd20178,15'd20177,15'd20176,15'd20175,15'd20174,15'd20173,15'd20172,15'd20171,15'd20170,15'd20169,15'd20168,15'd20167,15'd20166,15'd20165,15'd20164,15'd20163,15'd20162,15'd20161,15'd20160,
15'd19919,15'd19918,15'd19917,15'd19916,15'd19915,15'd19914,15'd19913,15'd19912,15'd19911,15'd19910,15'd19909,15'd19908,15'd19907,15'd19906,15'd19905,15'd19904,15'd19903,15'd19902,15'd19901,15'd19900,15'd19899,15'd19898,15'd19897,15'd19896,15'd19895,15'd19894,15'd19893,15'd19892,15'd19891,15'd19890,15'd19889,15'd19888,15'd19887,15'd19886,15'd19885,15'd19884,15'd19883,15'd19882,15'd19881,15'd19880,15'd19879,15'd19878,15'd19877,15'd19876,15'd19875,15'd19874,15'd19873,15'd19872,15'd19871,15'd19870,15'd19869,15'd19868,15'd19867,15'd19866,15'd19865,15'd19864,15'd19863,15'd19862,15'd19861,15'd19860,15'd19859,15'd19858,15'd19857,15'd19856,15'd19855,15'd19854,15'd19853,15'd19852,15'd19851,15'd19850,15'd19849,15'd19848,15'd19847,15'd19846,15'd19845,15'd19844,15'd19843,15'd19842,15'd19841,15'd19840,
15'd19599,15'd19598,15'd19597,15'd19596,15'd19595,15'd19594,15'd19593,15'd19592,15'd19591,15'd19590,15'd19589,15'd19588,15'd19587,15'd19586,15'd19585,15'd19584,15'd19583,15'd19582,15'd19581,15'd19580,15'd19579,15'd19578,15'd19577,15'd19576,15'd19575,15'd19574,15'd19573,15'd19572,15'd19571,15'd19570,15'd19569,15'd19568,15'd19567,15'd19566,15'd19565,15'd19564,15'd19563,15'd19562,15'd19561,15'd19560,15'd19559,15'd19558,15'd19557,15'd19556,15'd19555,15'd19554,15'd19553,15'd19552,15'd19551,15'd19550,15'd19549,15'd19548,15'd19547,15'd19546,15'd19545,15'd19544,15'd19543,15'd19542,15'd19541,15'd19540,15'd19539,15'd19538,15'd19537,15'd19536,15'd19535,15'd19534,15'd19533,15'd19532,15'd19531,15'd19530,15'd19529,15'd19528,15'd19527,15'd19526,15'd19525,15'd19524,15'd19523,15'd19522,15'd19521,15'd19520,
15'd19279,15'd19278,15'd19277,15'd19276,15'd19275,15'd19274,15'd19273,15'd19272,15'd19271,15'd19270,15'd19269,15'd19268,15'd19267,15'd19266,15'd19265,15'd19264,15'd19263,15'd19262,15'd19261,15'd19260,15'd19259,15'd19258,15'd19257,15'd19256,15'd19255,15'd19254,15'd19253,15'd19252,15'd19251,15'd19250,15'd19249,15'd19248,15'd19247,15'd19246,15'd19245,15'd19244,15'd19243,15'd19242,15'd19241,15'd19240,15'd19239,15'd19238,15'd19237,15'd19236,15'd19235,15'd19234,15'd19233,15'd19232,15'd19231,15'd19230,15'd19229,15'd19228,15'd19227,15'd19226,15'd19225,15'd19224,15'd19223,15'd19222,15'd19221,15'd19220,15'd19219,15'd19218,15'd19217,15'd19216,15'd19215,15'd19214,15'd19213,15'd19212,15'd19211,15'd19210,15'd19209,15'd19208,15'd19207,15'd19206,15'd19205,15'd19204,15'd19203,15'd19202,15'd19201,15'd19200,
15'd18959,15'd18958,15'd18957,15'd18956,15'd18955,15'd18954,15'd18953,15'd18952,15'd18951,15'd18950,15'd18949,15'd18948,15'd18947,15'd18946,15'd18945,15'd18944,15'd18943,15'd18942,15'd18941,15'd18940,15'd18939,15'd18938,15'd18937,15'd18936,15'd18935,15'd18934,15'd18933,15'd18932,15'd18931,15'd18930,15'd18929,15'd18928,15'd18927,15'd18926,15'd18925,15'd18924,15'd18923,15'd18922,15'd18921,15'd18920,15'd18919,15'd18918,15'd18917,15'd18916,15'd18915,15'd18914,15'd18913,15'd18912,15'd18911,15'd18910,15'd18909,15'd18908,15'd18907,15'd18906,15'd18905,15'd18904,15'd18903,15'd18902,15'd18901,15'd18900,15'd18899,15'd18898,15'd18897,15'd18896,15'd18895,15'd18894,15'd18893,15'd18892,15'd18891,15'd18890,15'd18889,15'd18888,15'd18887,15'd18886,15'd18885,15'd18884,15'd18883,15'd18882,15'd18881,15'd18880,
15'd18639,15'd18638,15'd18637,15'd18636,15'd18635,15'd18634,15'd18633,15'd18632,15'd18631,15'd18630,15'd18629,15'd18628,15'd18627,15'd18626,15'd18625,15'd18624,15'd18623,15'd18622,15'd18621,15'd18620,15'd18619,15'd18618,15'd18617,15'd18616,15'd18615,15'd18614,15'd18613,15'd18612,15'd18611,15'd18610,15'd18609,15'd18608,15'd18607,15'd18606,15'd18605,15'd18604,15'd18603,15'd18602,15'd18601,15'd18600,15'd18599,15'd18598,15'd18597,15'd18596,15'd18595,15'd18594,15'd18593,15'd18592,15'd18591,15'd18590,15'd18589,15'd18588,15'd18587,15'd18586,15'd18585,15'd18584,15'd18583,15'd18582,15'd18581,15'd18580,15'd18579,15'd18578,15'd18577,15'd18576,15'd18575,15'd18574,15'd18573,15'd18572,15'd18571,15'd18570,15'd18569,15'd18568,15'd18567,15'd18566,15'd18565,15'd18564,15'd18563,15'd18562,15'd18561,15'd18560,
15'd18319,15'd18318,15'd18317,15'd18316,15'd18315,15'd18314,15'd18313,15'd18312,15'd18311,15'd18310,15'd18309,15'd18308,15'd18307,15'd18306,15'd18305,15'd18304,15'd18303,15'd18302,15'd18301,15'd18300,15'd18299,15'd18298,15'd18297,15'd18296,15'd18295,15'd18294,15'd18293,15'd18292,15'd18291,15'd18290,15'd18289,15'd18288,15'd18287,15'd18286,15'd18285,15'd18284,15'd18283,15'd18282,15'd18281,15'd18280,15'd18279,15'd18278,15'd18277,15'd18276,15'd18275,15'd18274,15'd18273,15'd18272,15'd18271,15'd18270,15'd18269,15'd18268,15'd18267,15'd18266,15'd18265,15'd18264,15'd18263,15'd18262,15'd18261,15'd18260,15'd18259,15'd18258,15'd18257,15'd18256,15'd18255,15'd18254,15'd18253,15'd18252,15'd18251,15'd18250,15'd18249,15'd18248,15'd18247,15'd18246,15'd18245,15'd18244,15'd18243,15'd18242,15'd18241,15'd18240,
15'd17999,15'd17998,15'd17997,15'd17996,15'd17995,15'd17994,15'd17993,15'd17992,15'd17991,15'd17990,15'd17989,15'd17988,15'd17987,15'd17986,15'd17985,15'd17984,15'd17983,15'd17982,15'd17981,15'd17980,15'd17979,15'd17978,15'd17977,15'd17976,15'd17975,15'd17974,15'd17973,15'd17972,15'd17971,15'd17970,15'd17969,15'd17968,15'd17967,15'd17966,15'd17965,15'd17964,15'd17963,15'd17962,15'd17961,15'd17960,15'd17959,15'd17958,15'd17957,15'd17956,15'd17955,15'd17954,15'd17953,15'd17952,15'd17951,15'd17950,15'd17949,15'd17948,15'd17947,15'd17946,15'd17945,15'd17944,15'd17943,15'd17942,15'd17941,15'd17940,15'd17939,15'd17938,15'd17937,15'd17936,15'd17935,15'd17934,15'd17933,15'd17932,15'd17931,15'd17930,15'd17929,15'd17928,15'd17927,15'd17926,15'd17925,15'd17924,15'd17923,15'd17922,15'd17921,15'd17920,
15'd17679,15'd17678,15'd17677,15'd17676,15'd17675,15'd17674,15'd17673,15'd17672,15'd17671,15'd17670,15'd17669,15'd17668,15'd17667,15'd17666,15'd17665,15'd17664,15'd17663,15'd17662,15'd17661,15'd17660,15'd17659,15'd17658,15'd17657,15'd17656,15'd17655,15'd17654,15'd17653,15'd17652,15'd17651,15'd17650,15'd17649,15'd17648,15'd17647,15'd17646,15'd17645,15'd17644,15'd17643,15'd17642,15'd17641,15'd17640,15'd17639,15'd17638,15'd17637,15'd17636,15'd17635,15'd17634,15'd17633,15'd17632,15'd17631,15'd17630,15'd17629,15'd17628,15'd17627,15'd17626,15'd17625,15'd17624,15'd17623,15'd17622,15'd17621,15'd17620,15'd17619,15'd17618,15'd17617,15'd17616,15'd17615,15'd17614,15'd17613,15'd17612,15'd17611,15'd17610,15'd17609,15'd17608,15'd17607,15'd17606,15'd17605,15'd17604,15'd17603,15'd17602,15'd17601,15'd17600,
15'd17359,15'd17358,15'd17357,15'd17356,15'd17355,15'd17354,15'd17353,15'd17352,15'd17351,15'd17350,15'd17349,15'd17348,15'd17347,15'd17346,15'd17345,15'd17344,15'd17343,15'd17342,15'd17341,15'd17340,15'd17339,15'd17338,15'd17337,15'd17336,15'd17335,15'd17334,15'd17333,15'd17332,15'd17331,15'd17330,15'd17329,15'd17328,15'd17327,15'd17326,15'd17325,15'd17324,15'd17323,15'd17322,15'd17321,15'd17320,15'd17319,15'd17318,15'd17317,15'd17316,15'd17315,15'd17314,15'd17313,15'd17312,15'd17311,15'd17310,15'd17309,15'd17308,15'd17307,15'd17306,15'd17305,15'd17304,15'd17303,15'd17302,15'd17301,15'd17300,15'd17299,15'd17298,15'd17297,15'd17296,15'd17295,15'd17294,15'd17293,15'd17292,15'd17291,15'd17290,15'd17289,15'd17288,15'd17287,15'd17286,15'd17285,15'd17284,15'd17283,15'd17282,15'd17281,15'd17280,
15'd17039,15'd17038,15'd17037,15'd17036,15'd17035,15'd17034,15'd17033,15'd17032,15'd17031,15'd17030,15'd17029,15'd17028,15'd17027,15'd17026,15'd17025,15'd17024,15'd17023,15'd17022,15'd17021,15'd17020,15'd17019,15'd17018,15'd17017,15'd17016,15'd17015,15'd17014,15'd17013,15'd17012,15'd17011,15'd17010,15'd17009,15'd17008,15'd17007,15'd17006,15'd17005,15'd17004,15'd17003,15'd17002,15'd17001,15'd17000,15'd16999,15'd16998,15'd16997,15'd16996,15'd16995,15'd16994,15'd16993,15'd16992,15'd16991,15'd16990,15'd16989,15'd16988,15'd16987,15'd16986,15'd16985,15'd16984,15'd16983,15'd16982,15'd16981,15'd16980,15'd16979,15'd16978,15'd16977,15'd16976,15'd16975,15'd16974,15'd16973,15'd16972,15'd16971,15'd16970,15'd16969,15'd16968,15'd16967,15'd16966,15'd16965,15'd16964,15'd16963,15'd16962,15'd16961,15'd16960,
15'd16719,15'd16718,15'd16717,15'd16716,15'd16715,15'd16714,15'd16713,15'd16712,15'd16711,15'd16710,15'd16709,15'd16708,15'd16707,15'd16706,15'd16705,15'd16704,15'd16703,15'd16702,15'd16701,15'd16700,15'd16699,15'd16698,15'd16697,15'd16696,15'd16695,15'd16694,15'd16693,15'd16692,15'd16691,15'd16690,15'd16689,15'd16688,15'd16687,15'd16686,15'd16685,15'd16684,15'd16683,15'd16682,15'd16681,15'd16680,15'd16679,15'd16678,15'd16677,15'd16676,15'd16675,15'd16674,15'd16673,15'd16672,15'd16671,15'd16670,15'd16669,15'd16668,15'd16667,15'd16666,15'd16665,15'd16664,15'd16663,15'd16662,15'd16661,15'd16660,15'd16659,15'd16658,15'd16657,15'd16656,15'd16655,15'd16654,15'd16653,15'd16652,15'd16651,15'd16650,15'd16649,15'd16648,15'd16647,15'd16646,15'd16645,15'd16644,15'd16643,15'd16642,15'd16641,15'd16640,
15'd16399,15'd16398,15'd16397,15'd16396,15'd16395,15'd16394,15'd16393,15'd16392,15'd16391,15'd16390,15'd16389,15'd16388,15'd16387,15'd16386,15'd16385,15'd16384,15'd16383,15'd16382,15'd16381,15'd16380,15'd16379,15'd16378,15'd16377,15'd16376,15'd16375,15'd16374,15'd16373,15'd16372,15'd16371,15'd16370,15'd16369,15'd16368,15'd16367,15'd16366,15'd16365,15'd16364,15'd16363,15'd16362,15'd16361,15'd16360,15'd16359,15'd16358,15'd16357,15'd16356,15'd16355,15'd16354,15'd16353,15'd16352,15'd16351,15'd16350,15'd16349,15'd16348,15'd16347,15'd16346,15'd16345,15'd16344,15'd16343,15'd16342,15'd16341,15'd16340,15'd16339,15'd16338,15'd16337,15'd16336,15'd16335,15'd16334,15'd16333,15'd16332,15'd16331,15'd16330,15'd16329,15'd16328,15'd16327,15'd16326,15'd16325,15'd16324,15'd16323,15'd16322,15'd16321,15'd16320,
15'd16079,15'd16078,15'd16077,15'd16076,15'd16075,15'd16074,15'd16073,15'd16072,15'd16071,15'd16070,15'd16069,15'd16068,15'd16067,15'd16066,15'd16065,15'd16064,15'd16063,15'd16062,15'd16061,15'd16060,15'd16059,15'd16058,15'd16057,15'd16056,15'd16055,15'd16054,15'd16053,15'd16052,15'd16051,15'd16050,15'd16049,15'd16048,15'd16047,15'd16046,15'd16045,15'd16044,15'd16043,15'd16042,15'd16041,15'd16040,15'd16039,15'd16038,15'd16037,15'd16036,15'd16035,15'd16034,15'd16033,15'd16032,15'd16031,15'd16030,15'd16029,15'd16028,15'd16027,15'd16026,15'd16025,15'd16024,15'd16023,15'd16022,15'd16021,15'd16020,15'd16019,15'd16018,15'd16017,15'd16016,15'd16015,15'd16014,15'd16013,15'd16012,15'd16011,15'd16010,15'd16009,15'd16008,15'd16007,15'd16006,15'd16005,15'd16004,15'd16003,15'd16002,15'd16001,15'd16000,
15'd15759,15'd15758,15'd15757,15'd15756,15'd15755,15'd15754,15'd15753,15'd15752,15'd15751,15'd15750,15'd15749,15'd15748,15'd15747,15'd15746,15'd15745,15'd15744,15'd15743,15'd15742,15'd15741,15'd15740,15'd15739,15'd15738,15'd15737,15'd15736,15'd15735,15'd15734,15'd15733,15'd15732,15'd15731,15'd15730,15'd15729,15'd15728,15'd15727,15'd15726,15'd15725,15'd15724,15'd15723,15'd15722,15'd15721,15'd15720,15'd15719,15'd15718,15'd15717,15'd15716,15'd15715,15'd15714,15'd15713,15'd15712,15'd15711,15'd15710,15'd15709,15'd15708,15'd15707,15'd15706,15'd15705,15'd15704,15'd15703,15'd15702,15'd15701,15'd15700,15'd15699,15'd15698,15'd15697,15'd15696,15'd15695,15'd15694,15'd15693,15'd15692,15'd15691,15'd15690,15'd15689,15'd15688,15'd15687,15'd15686,15'd15685,15'd15684,15'd15683,15'd15682,15'd15681,15'd15680,
15'd15439,15'd15438,15'd15437,15'd15436,15'd15435,15'd15434,15'd15433,15'd15432,15'd15431,15'd15430,15'd15429,15'd15428,15'd15427,15'd15426,15'd15425,15'd15424,15'd15423,15'd15422,15'd15421,15'd15420,15'd15419,15'd15418,15'd15417,15'd15416,15'd15415,15'd15414,15'd15413,15'd15412,15'd15411,15'd15410,15'd15409,15'd15408,15'd15407,15'd15406,15'd15405,15'd15404,15'd15403,15'd15402,15'd15401,15'd15400,15'd15399,15'd15398,15'd15397,15'd15396,15'd15395,15'd15394,15'd15393,15'd15392,15'd15391,15'd15390,15'd15389,15'd15388,15'd15387,15'd15386,15'd15385,15'd15384,15'd15383,15'd15382,15'd15381,15'd15380,15'd15379,15'd15378,15'd15377,15'd15376,15'd15375,15'd15374,15'd15373,15'd15372,15'd15371,15'd15370,15'd15369,15'd15368,15'd15367,15'd15366,15'd15365,15'd15364,15'd15363,15'd15362,15'd15361,15'd15360,
15'd15119,15'd15118,15'd15117,15'd15116,15'd15115,15'd15114,15'd15113,15'd15112,15'd15111,15'd15110,15'd15109,15'd15108,15'd15107,15'd15106,15'd15105,15'd15104,15'd15103,15'd15102,15'd15101,15'd15100,15'd15099,15'd15098,15'd15097,15'd15096,15'd15095,15'd15094,15'd15093,15'd15092,15'd15091,15'd15090,15'd15089,15'd15088,15'd15087,15'd15086,15'd15085,15'd15084,15'd15083,15'd15082,15'd15081,15'd15080,15'd15079,15'd15078,15'd15077,15'd15076,15'd15075,15'd15074,15'd15073,15'd15072,15'd15071,15'd15070,15'd15069,15'd15068,15'd15067,15'd15066,15'd15065,15'd15064,15'd15063,15'd15062,15'd15061,15'd15060,15'd15059,15'd15058,15'd15057,15'd15056,15'd15055,15'd15054,15'd15053,15'd15052,15'd15051,15'd15050,15'd15049,15'd15048,15'd15047,15'd15046,15'd15045,15'd15044,15'd15043,15'd15042,15'd15041,15'd15040,
15'd14799,15'd14798,15'd14797,15'd14796,15'd14795,15'd14794,15'd14793,15'd14792,15'd14791,15'd14790,15'd14789,15'd14788,15'd14787,15'd14786,15'd14785,15'd14784,15'd14783,15'd14782,15'd14781,15'd14780,15'd14779,15'd14778,15'd14777,15'd14776,15'd14775,15'd14774,15'd14773,15'd14772,15'd14771,15'd14770,15'd14769,15'd14768,15'd14767,15'd14766,15'd14765,15'd14764,15'd14763,15'd14762,15'd14761,15'd14760,15'd14759,15'd14758,15'd14757,15'd14756,15'd14755,15'd14754,15'd14753,15'd14752,15'd14751,15'd14750,15'd14749,15'd14748,15'd14747,15'd14746,15'd14745,15'd14744,15'd14743,15'd14742,15'd14741,15'd14740,15'd14739,15'd14738,15'd14737,15'd14736,15'd14735,15'd14734,15'd14733,15'd14732,15'd14731,15'd14730,15'd14729,15'd14728,15'd14727,15'd14726,15'd14725,15'd14724,15'd14723,15'd14722,15'd14721,15'd14720,
15'd14479,15'd14478,15'd14477,15'd14476,15'd14475,15'd14474,15'd14473,15'd14472,15'd14471,15'd14470,15'd14469,15'd14468,15'd14467,15'd14466,15'd14465,15'd14464,15'd14463,15'd14462,15'd14461,15'd14460,15'd14459,15'd14458,15'd14457,15'd14456,15'd14455,15'd14454,15'd14453,15'd14452,15'd14451,15'd14450,15'd14449,15'd14448,15'd14447,15'd14446,15'd14445,15'd14444,15'd14443,15'd14442,15'd14441,15'd14440,15'd14439,15'd14438,15'd14437,15'd14436,15'd14435,15'd14434,15'd14433,15'd14432,15'd14431,15'd14430,15'd14429,15'd14428,15'd14427,15'd14426,15'd14425,15'd14424,15'd14423,15'd14422,15'd14421,15'd14420,15'd14419,15'd14418,15'd14417,15'd14416,15'd14415,15'd14414,15'd14413,15'd14412,15'd14411,15'd14410,15'd14409,15'd14408,15'd14407,15'd14406,15'd14405,15'd14404,15'd14403,15'd14402,15'd14401,15'd14400,
15'd14159,15'd14158,15'd14157,15'd14156,15'd14155,15'd14154,15'd14153,15'd14152,15'd14151,15'd14150,15'd14149,15'd14148,15'd14147,15'd14146,15'd14145,15'd14144,15'd14143,15'd14142,15'd14141,15'd14140,15'd14139,15'd14138,15'd14137,15'd14136,15'd14135,15'd14134,15'd14133,15'd14132,15'd14131,15'd14130,15'd14129,15'd14128,15'd14127,15'd14126,15'd14125,15'd14124,15'd14123,15'd14122,15'd14121,15'd14120,15'd14119,15'd14118,15'd14117,15'd14116,15'd14115,15'd14114,15'd14113,15'd14112,15'd14111,15'd14110,15'd14109,15'd14108,15'd14107,15'd14106,15'd14105,15'd14104,15'd14103,15'd14102,15'd14101,15'd14100,15'd14099,15'd14098,15'd14097,15'd14096,15'd14095,15'd14094,15'd14093,15'd14092,15'd14091,15'd14090,15'd14089,15'd14088,15'd14087,15'd14086,15'd14085,15'd14084,15'd14083,15'd14082,15'd14081,15'd14080,
15'd13839,15'd13838,15'd13837,15'd13836,15'd13835,15'd13834,15'd13833,15'd13832,15'd13831,15'd13830,15'd13829,15'd13828,15'd13827,15'd13826,15'd13825,15'd13824,15'd13823,15'd13822,15'd13821,15'd13820,15'd13819,15'd13818,15'd13817,15'd13816,15'd13815,15'd13814,15'd13813,15'd13812,15'd13811,15'd13810,15'd13809,15'd13808,15'd13807,15'd13806,15'd13805,15'd13804,15'd13803,15'd13802,15'd13801,15'd13800,15'd13799,15'd13798,15'd13797,15'd13796,15'd13795,15'd13794,15'd13793,15'd13792,15'd13791,15'd13790,15'd13789,15'd13788,15'd13787,15'd13786,15'd13785,15'd13784,15'd13783,15'd13782,15'd13781,15'd13780,15'd13779,15'd13778,15'd13777,15'd13776,15'd13775,15'd13774,15'd13773,15'd13772,15'd13771,15'd13770,15'd13769,15'd13768,15'd13767,15'd13766,15'd13765,15'd13764,15'd13763,15'd13762,15'd13761,15'd13760,
15'd13519,15'd13518,15'd13517,15'd13516,15'd13515,15'd13514,15'd13513,15'd13512,15'd13511,15'd13510,15'd13509,15'd13508,15'd13507,15'd13506,15'd13505,15'd13504,15'd13503,15'd13502,15'd13501,15'd13500,15'd13499,15'd13498,15'd13497,15'd13496,15'd13495,15'd13494,15'd13493,15'd13492,15'd13491,15'd13490,15'd13489,15'd13488,15'd13487,15'd13486,15'd13485,15'd13484,15'd13483,15'd13482,15'd13481,15'd13480,15'd13479,15'd13478,15'd13477,15'd13476,15'd13475,15'd13474,15'd13473,15'd13472,15'd13471,15'd13470,15'd13469,15'd13468,15'd13467,15'd13466,15'd13465,15'd13464,15'd13463,15'd13462,15'd13461,15'd13460,15'd13459,15'd13458,15'd13457,15'd13456,15'd13455,15'd13454,15'd13453,15'd13452,15'd13451,15'd13450,15'd13449,15'd13448,15'd13447,15'd13446,15'd13445,15'd13444,15'd13443,15'd13442,15'd13441,15'd13440,
15'd13199,15'd13198,15'd13197,15'd13196,15'd13195,15'd13194,15'd13193,15'd13192,15'd13191,15'd13190,15'd13189,15'd13188,15'd13187,15'd13186,15'd13185,15'd13184,15'd13183,15'd13182,15'd13181,15'd13180,15'd13179,15'd13178,15'd13177,15'd13176,15'd13175,15'd13174,15'd13173,15'd13172,15'd13171,15'd13170,15'd13169,15'd13168,15'd13167,15'd13166,15'd13165,15'd13164,15'd13163,15'd13162,15'd13161,15'd13160,15'd13159,15'd13158,15'd13157,15'd13156,15'd13155,15'd13154,15'd13153,15'd13152,15'd13151,15'd13150,15'd13149,15'd13148,15'd13147,15'd13146,15'd13145,15'd13144,15'd13143,15'd13142,15'd13141,15'd13140,15'd13139,15'd13138,15'd13137,15'd13136,15'd13135,15'd13134,15'd13133,15'd13132,15'd13131,15'd13130,15'd13129,15'd13128,15'd13127,15'd13126,15'd13125,15'd13124,15'd13123,15'd13122,15'd13121,15'd13120,
15'd12879,15'd12878,15'd12877,15'd12876,15'd12875,15'd12874,15'd12873,15'd12872,15'd12871,15'd12870,15'd12869,15'd12868,15'd12867,15'd12866,15'd12865,15'd12864,15'd12863,15'd12862,15'd12861,15'd12860,15'd12859,15'd12858,15'd12857,15'd12856,15'd12855,15'd12854,15'd12853,15'd12852,15'd12851,15'd12850,15'd12849,15'd12848,15'd12847,15'd12846,15'd12845,15'd12844,15'd12843,15'd12842,15'd12841,15'd12840,15'd12839,15'd12838,15'd12837,15'd12836,15'd12835,15'd12834,15'd12833,15'd12832,15'd12831,15'd12830,15'd12829,15'd12828,15'd12827,15'd12826,15'd12825,15'd12824,15'd12823,15'd12822,15'd12821,15'd12820,15'd12819,15'd12818,15'd12817,15'd12816,15'd12815,15'd12814,15'd12813,15'd12812,15'd12811,15'd12810,15'd12809,15'd12808,15'd12807,15'd12806,15'd12805,15'd12804,15'd12803,15'd12802,15'd12801,15'd12800,
15'd12559,15'd12558,15'd12557,15'd12556,15'd12555,15'd12554,15'd12553,15'd12552,15'd12551,15'd12550,15'd12549,15'd12548,15'd12547,15'd12546,15'd12545,15'd12544,15'd12543,15'd12542,15'd12541,15'd12540,15'd12539,15'd12538,15'd12537,15'd12536,15'd12535,15'd12534,15'd12533,15'd12532,15'd12531,15'd12530,15'd12529,15'd12528,15'd12527,15'd12526,15'd12525,15'd12524,15'd12523,15'd12522,15'd12521,15'd12520,15'd12519,15'd12518,15'd12517,15'd12516,15'd12515,15'd12514,15'd12513,15'd12512,15'd12511,15'd12510,15'd12509,15'd12508,15'd12507,15'd12506,15'd12505,15'd12504,15'd12503,15'd12502,15'd12501,15'd12500,15'd12499,15'd12498,15'd12497,15'd12496,15'd12495,15'd12494,15'd12493,15'd12492,15'd12491,15'd12490,15'd12489,15'd12488,15'd12487,15'd12486,15'd12485,15'd12484,15'd12483,15'd12482,15'd12481,15'd12480,
15'd12239,15'd12238,15'd12237,15'd12236,15'd12235,15'd12234,15'd12233,15'd12232,15'd12231,15'd12230,15'd12229,15'd12228,15'd12227,15'd12226,15'd12225,15'd12224,15'd12223,15'd12222,15'd12221,15'd12220,15'd12219,15'd12218,15'd12217,15'd12216,15'd12215,15'd12214,15'd12213,15'd12212,15'd12211,15'd12210,15'd12209,15'd12208,15'd12207,15'd12206,15'd12205,15'd12204,15'd12203,15'd12202,15'd12201,15'd12200,15'd12199,15'd12198,15'd12197,15'd12196,15'd12195,15'd12194,15'd12193,15'd12192,15'd12191,15'd12190,15'd12189,15'd12188,15'd12187,15'd12186,15'd12185,15'd12184,15'd12183,15'd12182,15'd12181,15'd12180,15'd12179,15'd12178,15'd12177,15'd12176,15'd12175,15'd12174,15'd12173,15'd12172,15'd12171,15'd12170,15'd12169,15'd12168,15'd12167,15'd12166,15'd12165,15'd12164,15'd12163,15'd12162,15'd12161,15'd12160,
15'd11919,15'd11918,15'd11917,15'd11916,15'd11915,15'd11914,15'd11913,15'd11912,15'd11911,15'd11910,15'd11909,15'd11908,15'd11907,15'd11906,15'd11905,15'd11904,15'd11903,15'd11902,15'd11901,15'd11900,15'd11899,15'd11898,15'd11897,15'd11896,15'd11895,15'd11894,15'd11893,15'd11892,15'd11891,15'd11890,15'd11889,15'd11888,15'd11887,15'd11886,15'd11885,15'd11884,15'd11883,15'd11882,15'd11881,15'd11880,15'd11879,15'd11878,15'd11877,15'd11876,15'd11875,15'd11874,15'd11873,15'd11872,15'd11871,15'd11870,15'd11869,15'd11868,15'd11867,15'd11866,15'd11865,15'd11864,15'd11863,15'd11862,15'd11861,15'd11860,15'd11859,15'd11858,15'd11857,15'd11856,15'd11855,15'd11854,15'd11853,15'd11852,15'd11851,15'd11850,15'd11849,15'd11848,15'd11847,15'd11846,15'd11845,15'd11844,15'd11843,15'd11842,15'd11841,15'd11840,
15'd11599,15'd11598,15'd11597,15'd11596,15'd11595,15'd11594,15'd11593,15'd11592,15'd11591,15'd11590,15'd11589,15'd11588,15'd11587,15'd11586,15'd11585,15'd11584,15'd11583,15'd11582,15'd11581,15'd11580,15'd11579,15'd11578,15'd11577,15'd11576,15'd11575,15'd11574,15'd11573,15'd11572,15'd11571,15'd11570,15'd11569,15'd11568,15'd11567,15'd11566,15'd11565,15'd11564,15'd11563,15'd11562,15'd11561,15'd11560,15'd11559,15'd11558,15'd11557,15'd11556,15'd11555,15'd11554,15'd11553,15'd11552,15'd11551,15'd11550,15'd11549,15'd11548,15'd11547,15'd11546,15'd11545,15'd11544,15'd11543,15'd11542,15'd11541,15'd11540,15'd11539,15'd11538,15'd11537,15'd11536,15'd11535,15'd11534,15'd11533,15'd11532,15'd11531,15'd11530,15'd11529,15'd11528,15'd11527,15'd11526,15'd11525,15'd11524,15'd11523,15'd11522,15'd11521,15'd11520,
15'd11279,15'd11278,15'd11277,15'd11276,15'd11275,15'd11274,15'd11273,15'd11272,15'd11271,15'd11270,15'd11269,15'd11268,15'd11267,15'd11266,15'd11265,15'd11264,15'd11263,15'd11262,15'd11261,15'd11260,15'd11259,15'd11258,15'd11257,15'd11256,15'd11255,15'd11254,15'd11253,15'd11252,15'd11251,15'd11250,15'd11249,15'd11248,15'd11247,15'd11246,15'd11245,15'd11244,15'd11243,15'd11242,15'd11241,15'd11240,15'd11239,15'd11238,15'd11237,15'd11236,15'd11235,15'd11234,15'd11233,15'd11232,15'd11231,15'd11230,15'd11229,15'd11228,15'd11227,15'd11226,15'd11225,15'd11224,15'd11223,15'd11222,15'd11221,15'd11220,15'd11219,15'd11218,15'd11217,15'd11216,15'd11215,15'd11214,15'd11213,15'd11212,15'd11211,15'd11210,15'd11209,15'd11208,15'd11207,15'd11206,15'd11205,15'd11204,15'd11203,15'd11202,15'd11201,15'd11200,
15'd10959,15'd10958,15'd10957,15'd10956,15'd10955,15'd10954,15'd10953,15'd10952,15'd10951,15'd10950,15'd10949,15'd10948,15'd10947,15'd10946,15'd10945,15'd10944,15'd10943,15'd10942,15'd10941,15'd10940,15'd10939,15'd10938,15'd10937,15'd10936,15'd10935,15'd10934,15'd10933,15'd10932,15'd10931,15'd10930,15'd10929,15'd10928,15'd10927,15'd10926,15'd10925,15'd10924,15'd10923,15'd10922,15'd10921,15'd10920,15'd10919,15'd10918,15'd10917,15'd10916,15'd10915,15'd10914,15'd10913,15'd10912,15'd10911,15'd10910,15'd10909,15'd10908,15'd10907,15'd10906,15'd10905,15'd10904,15'd10903,15'd10902,15'd10901,15'd10900,15'd10899,15'd10898,15'd10897,15'd10896,15'd10895,15'd10894,15'd10893,15'd10892,15'd10891,15'd10890,15'd10889,15'd10888,15'd10887,15'd10886,15'd10885,15'd10884,15'd10883,15'd10882,15'd10881,15'd10880,
15'd10639,15'd10638,15'd10637,15'd10636,15'd10635,15'd10634,15'd10633,15'd10632,15'd10631,15'd10630,15'd10629,15'd10628,15'd10627,15'd10626,15'd10625,15'd10624,15'd10623,15'd10622,15'd10621,15'd10620,15'd10619,15'd10618,15'd10617,15'd10616,15'd10615,15'd10614,15'd10613,15'd10612,15'd10611,15'd10610,15'd10609,15'd10608,15'd10607,15'd10606,15'd10605,15'd10604,15'd10603,15'd10602,15'd10601,15'd10600,15'd10599,15'd10598,15'd10597,15'd10596,15'd10595,15'd10594,15'd10593,15'd10592,15'd10591,15'd10590,15'd10589,15'd10588,15'd10587,15'd10586,15'd10585,15'd10584,15'd10583,15'd10582,15'd10581,15'd10580,15'd10579,15'd10578,15'd10577,15'd10576,15'd10575,15'd10574,15'd10573,15'd10572,15'd10571,15'd10570,15'd10569,15'd10568,15'd10567,15'd10566,15'd10565,15'd10564,15'd10563,15'd10562,15'd10561,15'd10560,
15'd10319,15'd10318,15'd10317,15'd10316,15'd10315,15'd10314,15'd10313,15'd10312,15'd10311,15'd10310,15'd10309,15'd10308,15'd10307,15'd10306,15'd10305,15'd10304,15'd10303,15'd10302,15'd10301,15'd10300,15'd10299,15'd10298,15'd10297,15'd10296,15'd10295,15'd10294,15'd10293,15'd10292,15'd10291,15'd10290,15'd10289,15'd10288,15'd10287,15'd10286,15'd10285,15'd10284,15'd10283,15'd10282,15'd10281,15'd10280,15'd10279,15'd10278,15'd10277,15'd10276,15'd10275,15'd10274,15'd10273,15'd10272,15'd10271,15'd10270,15'd10269,15'd10268,15'd10267,15'd10266,15'd10265,15'd10264,15'd10263,15'd10262,15'd10261,15'd10260,15'd10259,15'd10258,15'd10257,15'd10256,15'd10255,15'd10254,15'd10253,15'd10252,15'd10251,15'd10250,15'd10249,15'd10248,15'd10247,15'd10246,15'd10245,15'd10244,15'd10243,15'd10242,15'd10241,15'd10240,
15'd9999,15'd9998,15'd9997,15'd9996,15'd9995,15'd9994,15'd9993,15'd9992,15'd9991,15'd9990,15'd9989,15'd9988,15'd9987,15'd9986,15'd9985,15'd9984,15'd9983,15'd9982,15'd9981,15'd9980,15'd9979,15'd9978,15'd9977,15'd9976,15'd9975,15'd9974,15'd9973,15'd9972,15'd9971,15'd9970,15'd9969,15'd9968,15'd9967,15'd9966,15'd9965,15'd9964,15'd9963,15'd9962,15'd9961,15'd9960,15'd9959,15'd9958,15'd9957,15'd9956,15'd9955,15'd9954,15'd9953,15'd9952,15'd9951,15'd9950,15'd9949,15'd9948,15'd9947,15'd9946,15'd9945,15'd9944,15'd9943,15'd9942,15'd9941,15'd9940,15'd9939,15'd9938,15'd9937,15'd9936,15'd9935,15'd9934,15'd9933,15'd9932,15'd9931,15'd9930,15'd9929,15'd9928,15'd9927,15'd9926,15'd9925,15'd9924,15'd9923,15'd9922,15'd9921,15'd9920,
15'd9679,15'd9678,15'd9677,15'd9676,15'd9675,15'd9674,15'd9673,15'd9672,15'd9671,15'd9670,15'd9669,15'd9668,15'd9667,15'd9666,15'd9665,15'd9664,15'd9663,15'd9662,15'd9661,15'd9660,15'd9659,15'd9658,15'd9657,15'd9656,15'd9655,15'd9654,15'd9653,15'd9652,15'd9651,15'd9650,15'd9649,15'd9648,15'd9647,15'd9646,15'd9645,15'd9644,15'd9643,15'd9642,15'd9641,15'd9640,15'd9639,15'd9638,15'd9637,15'd9636,15'd9635,15'd9634,15'd9633,15'd9632,15'd9631,15'd9630,15'd9629,15'd9628,15'd9627,15'd9626,15'd9625,15'd9624,15'd9623,15'd9622,15'd9621,15'd9620,15'd9619,15'd9618,15'd9617,15'd9616,15'd9615,15'd9614,15'd9613,15'd9612,15'd9611,15'd9610,15'd9609,15'd9608,15'd9607,15'd9606,15'd9605,15'd9604,15'd9603,15'd9602,15'd9601,15'd9600,
15'd9359,15'd9358,15'd9357,15'd9356,15'd9355,15'd9354,15'd9353,15'd9352,15'd9351,15'd9350,15'd9349,15'd9348,15'd9347,15'd9346,15'd9345,15'd9344,15'd9343,15'd9342,15'd9341,15'd9340,15'd9339,15'd9338,15'd9337,15'd9336,15'd9335,15'd9334,15'd9333,15'd9332,15'd9331,15'd9330,15'd9329,15'd9328,15'd9327,15'd9326,15'd9325,15'd9324,15'd9323,15'd9322,15'd9321,15'd9320,15'd9319,15'd9318,15'd9317,15'd9316,15'd9315,15'd9314,15'd9313,15'd9312,15'd9311,15'd9310,15'd9309,15'd9308,15'd9307,15'd9306,15'd9305,15'd9304,15'd9303,15'd9302,15'd9301,15'd9300,15'd9299,15'd9298,15'd9297,15'd9296,15'd9295,15'd9294,15'd9293,15'd9292,15'd9291,15'd9290,15'd9289,15'd9288,15'd9287,15'd9286,15'd9285,15'd9284,15'd9283,15'd9282,15'd9281,15'd9280,
15'd9039,15'd9038,15'd9037,15'd9036,15'd9035,15'd9034,15'd9033,15'd9032,15'd9031,15'd9030,15'd9029,15'd9028,15'd9027,15'd9026,15'd9025,15'd9024,15'd9023,15'd9022,15'd9021,15'd9020,15'd9019,15'd9018,15'd9017,15'd9016,15'd9015,15'd9014,15'd9013,15'd9012,15'd9011,15'd9010,15'd9009,15'd9008,15'd9007,15'd9006,15'd9005,15'd9004,15'd9003,15'd9002,15'd9001,15'd9000,15'd8999,15'd8998,15'd8997,15'd8996,15'd8995,15'd8994,15'd8993,15'd8992,15'd8991,15'd8990,15'd8989,15'd8988,15'd8987,15'd8986,15'd8985,15'd8984,15'd8983,15'd8982,15'd8981,15'd8980,15'd8979,15'd8978,15'd8977,15'd8976,15'd8975,15'd8974,15'd8973,15'd8972,15'd8971,15'd8970,15'd8969,15'd8968,15'd8967,15'd8966,15'd8965,15'd8964,15'd8963,15'd8962,15'd8961,15'd8960,
15'd8719,15'd8718,15'd8717,15'd8716,15'd8715,15'd8714,15'd8713,15'd8712,15'd8711,15'd8710,15'd8709,15'd8708,15'd8707,15'd8706,15'd8705,15'd8704,15'd8703,15'd8702,15'd8701,15'd8700,15'd8699,15'd8698,15'd8697,15'd8696,15'd8695,15'd8694,15'd8693,15'd8692,15'd8691,15'd8690,15'd8689,15'd8688,15'd8687,15'd8686,15'd8685,15'd8684,15'd8683,15'd8682,15'd8681,15'd8680,15'd8679,15'd8678,15'd8677,15'd8676,15'd8675,15'd8674,15'd8673,15'd8672,15'd8671,15'd8670,15'd8669,15'd8668,15'd8667,15'd8666,15'd8665,15'd8664,15'd8663,15'd8662,15'd8661,15'd8660,15'd8659,15'd8658,15'd8657,15'd8656,15'd8655,15'd8654,15'd8653,15'd8652,15'd8651,15'd8650,15'd8649,15'd8648,15'd8647,15'd8646,15'd8645,15'd8644,15'd8643,15'd8642,15'd8641,15'd8640,
15'd8399,15'd8398,15'd8397,15'd8396,15'd8395,15'd8394,15'd8393,15'd8392,15'd8391,15'd8390,15'd8389,15'd8388,15'd8387,15'd8386,15'd8385,15'd8384,15'd8383,15'd8382,15'd8381,15'd8380,15'd8379,15'd8378,15'd8377,15'd8376,15'd8375,15'd8374,15'd8373,15'd8372,15'd8371,15'd8370,15'd8369,15'd8368,15'd8367,15'd8366,15'd8365,15'd8364,15'd8363,15'd8362,15'd8361,15'd8360,15'd8359,15'd8358,15'd8357,15'd8356,15'd8355,15'd8354,15'd8353,15'd8352,15'd8351,15'd8350,15'd8349,15'd8348,15'd8347,15'd8346,15'd8345,15'd8344,15'd8343,15'd8342,15'd8341,15'd8340,15'd8339,15'd8338,15'd8337,15'd8336,15'd8335,15'd8334,15'd8333,15'd8332,15'd8331,15'd8330,15'd8329,15'd8328,15'd8327,15'd8326,15'd8325,15'd8324,15'd8323,15'd8322,15'd8321,15'd8320,
15'd8079,15'd8078,15'd8077,15'd8076,15'd8075,15'd8074,15'd8073,15'd8072,15'd8071,15'd8070,15'd8069,15'd8068,15'd8067,15'd8066,15'd8065,15'd8064,15'd8063,15'd8062,15'd8061,15'd8060,15'd8059,15'd8058,15'd8057,15'd8056,15'd8055,15'd8054,15'd8053,15'd8052,15'd8051,15'd8050,15'd8049,15'd8048,15'd8047,15'd8046,15'd8045,15'd8044,15'd8043,15'd8042,15'd8041,15'd8040,15'd8039,15'd8038,15'd8037,15'd8036,15'd8035,15'd8034,15'd8033,15'd8032,15'd8031,15'd8030,15'd8029,15'd8028,15'd8027,15'd8026,15'd8025,15'd8024,15'd8023,15'd8022,15'd8021,15'd8020,15'd8019,15'd8018,15'd8017,15'd8016,15'd8015,15'd8014,15'd8013,15'd8012,15'd8011,15'd8010,15'd8009,15'd8008,15'd8007,15'd8006,15'd8005,15'd8004,15'd8003,15'd8002,15'd8001,15'd8000,
15'd7759,15'd7758,15'd7757,15'd7756,15'd7755,15'd7754,15'd7753,15'd7752,15'd7751,15'd7750,15'd7749,15'd7748,15'd7747,15'd7746,15'd7745,15'd7744,15'd7743,15'd7742,15'd7741,15'd7740,15'd7739,15'd7738,15'd7737,15'd7736,15'd7735,15'd7734,15'd7733,15'd7732,15'd7731,15'd7730,15'd7729,15'd7728,15'd7727,15'd7726,15'd7725,15'd7724,15'd7723,15'd7722,15'd7721,15'd7720,15'd7719,15'd7718,15'd7717,15'd7716,15'd7715,15'd7714,15'd7713,15'd7712,15'd7711,15'd7710,15'd7709,15'd7708,15'd7707,15'd7706,15'd7705,15'd7704,15'd7703,15'd7702,15'd7701,15'd7700,15'd7699,15'd7698,15'd7697,15'd7696,15'd7695,15'd7694,15'd7693,15'd7692,15'd7691,15'd7690,15'd7689,15'd7688,15'd7687,15'd7686,15'd7685,15'd7684,15'd7683,15'd7682,15'd7681,15'd7680,
15'd7439,15'd7438,15'd7437,15'd7436,15'd7435,15'd7434,15'd7433,15'd7432,15'd7431,15'd7430,15'd7429,15'd7428,15'd7427,15'd7426,15'd7425,15'd7424,15'd7423,15'd7422,15'd7421,15'd7420,15'd7419,15'd7418,15'd7417,15'd7416,15'd7415,15'd7414,15'd7413,15'd7412,15'd7411,15'd7410,15'd7409,15'd7408,15'd7407,15'd7406,15'd7405,15'd7404,15'd7403,15'd7402,15'd7401,15'd7400,15'd7399,15'd7398,15'd7397,15'd7396,15'd7395,15'd7394,15'd7393,15'd7392,15'd7391,15'd7390,15'd7389,15'd7388,15'd7387,15'd7386,15'd7385,15'd7384,15'd7383,15'd7382,15'd7381,15'd7380,15'd7379,15'd7378,15'd7377,15'd7376,15'd7375,15'd7374,15'd7373,15'd7372,15'd7371,15'd7370,15'd7369,15'd7368,15'd7367,15'd7366,15'd7365,15'd7364,15'd7363,15'd7362,15'd7361,15'd7360,
15'd7119,15'd7118,15'd7117,15'd7116,15'd7115,15'd7114,15'd7113,15'd7112,15'd7111,15'd7110,15'd7109,15'd7108,15'd7107,15'd7106,15'd7105,15'd7104,15'd7103,15'd7102,15'd7101,15'd7100,15'd7099,15'd7098,15'd7097,15'd7096,15'd7095,15'd7094,15'd7093,15'd7092,15'd7091,15'd7090,15'd7089,15'd7088,15'd7087,15'd7086,15'd7085,15'd7084,15'd7083,15'd7082,15'd7081,15'd7080,15'd7079,15'd7078,15'd7077,15'd7076,15'd7075,15'd7074,15'd7073,15'd7072,15'd7071,15'd7070,15'd7069,15'd7068,15'd7067,15'd7066,15'd7065,15'd7064,15'd7063,15'd7062,15'd7061,15'd7060,15'd7059,15'd7058,15'd7057,15'd7056,15'd7055,15'd7054,15'd7053,15'd7052,15'd7051,15'd7050,15'd7049,15'd7048,15'd7047,15'd7046,15'd7045,15'd7044,15'd7043,15'd7042,15'd7041,15'd7040,
15'd6799,15'd6798,15'd6797,15'd6796,15'd6795,15'd6794,15'd6793,15'd6792,15'd6791,15'd6790,15'd6789,15'd6788,15'd6787,15'd6786,15'd6785,15'd6784,15'd6783,15'd6782,15'd6781,15'd6780,15'd6779,15'd6778,15'd6777,15'd6776,15'd6775,15'd6774,15'd6773,15'd6772,15'd6771,15'd6770,15'd6769,15'd6768,15'd6767,15'd6766,15'd6765,15'd6764,15'd6763,15'd6762,15'd6761,15'd6760,15'd6759,15'd6758,15'd6757,15'd6756,15'd6755,15'd6754,15'd6753,15'd6752,15'd6751,15'd6750,15'd6749,15'd6748,15'd6747,15'd6746,15'd6745,15'd6744,15'd6743,15'd6742,15'd6741,15'd6740,15'd6739,15'd6738,15'd6737,15'd6736,15'd6735,15'd6734,15'd6733,15'd6732,15'd6731,15'd6730,15'd6729,15'd6728,15'd6727,15'd6726,15'd6725,15'd6724,15'd6723,15'd6722,15'd6721,15'd6720,
15'd6479,15'd6478,15'd6477,15'd6476,15'd6475,15'd6474,15'd6473,15'd6472,15'd6471,15'd6470,15'd6469,15'd6468,15'd6467,15'd6466,15'd6465,15'd6464,15'd6463,15'd6462,15'd6461,15'd6460,15'd6459,15'd6458,15'd6457,15'd6456,15'd6455,15'd6454,15'd6453,15'd6452,15'd6451,15'd6450,15'd6449,15'd6448,15'd6447,15'd6446,15'd6445,15'd6444,15'd6443,15'd6442,15'd6441,15'd6440,15'd6439,15'd6438,15'd6437,15'd6436,15'd6435,15'd6434,15'd6433,15'd6432,15'd6431,15'd6430,15'd6429,15'd6428,15'd6427,15'd6426,15'd6425,15'd6424,15'd6423,15'd6422,15'd6421,15'd6420,15'd6419,15'd6418,15'd6417,15'd6416,15'd6415,15'd6414,15'd6413,15'd6412,15'd6411,15'd6410,15'd6409,15'd6408,15'd6407,15'd6406,15'd6405,15'd6404,15'd6403,15'd6402,15'd6401,15'd6400,
15'd6159,15'd6158,15'd6157,15'd6156,15'd6155,15'd6154,15'd6153,15'd6152,15'd6151,15'd6150,15'd6149,15'd6148,15'd6147,15'd6146,15'd6145,15'd6144,15'd6143,15'd6142,15'd6141,15'd6140,15'd6139,15'd6138,15'd6137,15'd6136,15'd6135,15'd6134,15'd6133,15'd6132,15'd6131,15'd6130,15'd6129,15'd6128,15'd6127,15'd6126,15'd6125,15'd6124,15'd6123,15'd6122,15'd6121,15'd6120,15'd6119,15'd6118,15'd6117,15'd6116,15'd6115,15'd6114,15'd6113,15'd6112,15'd6111,15'd6110,15'd6109,15'd6108,15'd6107,15'd6106,15'd6105,15'd6104,15'd6103,15'd6102,15'd6101,15'd6100,15'd6099,15'd6098,15'd6097,15'd6096,15'd6095,15'd6094,15'd6093,15'd6092,15'd6091,15'd6090,15'd6089,15'd6088,15'd6087,15'd6086,15'd6085,15'd6084,15'd6083,15'd6082,15'd6081,15'd6080,
15'd5839,15'd5838,15'd5837,15'd5836,15'd5835,15'd5834,15'd5833,15'd5832,15'd5831,15'd5830,15'd5829,15'd5828,15'd5827,15'd5826,15'd5825,15'd5824,15'd5823,15'd5822,15'd5821,15'd5820,15'd5819,15'd5818,15'd5817,15'd5816,15'd5815,15'd5814,15'd5813,15'd5812,15'd5811,15'd5810,15'd5809,15'd5808,15'd5807,15'd5806,15'd5805,15'd5804,15'd5803,15'd5802,15'd5801,15'd5800,15'd5799,15'd5798,15'd5797,15'd5796,15'd5795,15'd5794,15'd5793,15'd5792,15'd5791,15'd5790,15'd5789,15'd5788,15'd5787,15'd5786,15'd5785,15'd5784,15'd5783,15'd5782,15'd5781,15'd5780,15'd5779,15'd5778,15'd5777,15'd5776,15'd5775,15'd5774,15'd5773,15'd5772,15'd5771,15'd5770,15'd5769,15'd5768,15'd5767,15'd5766,15'd5765,15'd5764,15'd5763,15'd5762,15'd5761,15'd5760,
15'd5519,15'd5518,15'd5517,15'd5516,15'd5515,15'd5514,15'd5513,15'd5512,15'd5511,15'd5510,15'd5509,15'd5508,15'd5507,15'd5506,15'd5505,15'd5504,15'd5503,15'd5502,15'd5501,15'd5500,15'd5499,15'd5498,15'd5497,15'd5496,15'd5495,15'd5494,15'd5493,15'd5492,15'd5491,15'd5490,15'd5489,15'd5488,15'd5487,15'd5486,15'd5485,15'd5484,15'd5483,15'd5482,15'd5481,15'd5480,15'd5479,15'd5478,15'd5477,15'd5476,15'd5475,15'd5474,15'd5473,15'd5472,15'd5471,15'd5470,15'd5469,15'd5468,15'd5467,15'd5466,15'd5465,15'd5464,15'd5463,15'd5462,15'd5461,15'd5460,15'd5459,15'd5458,15'd5457,15'd5456,15'd5455,15'd5454,15'd5453,15'd5452,15'd5451,15'd5450,15'd5449,15'd5448,15'd5447,15'd5446,15'd5445,15'd5444,15'd5443,15'd5442,15'd5441,15'd5440,
15'd5199,15'd5198,15'd5197,15'd5196,15'd5195,15'd5194,15'd5193,15'd5192,15'd5191,15'd5190,15'd5189,15'd5188,15'd5187,15'd5186,15'd5185,15'd5184,15'd5183,15'd5182,15'd5181,15'd5180,15'd5179,15'd5178,15'd5177,15'd5176,15'd5175,15'd5174,15'd5173,15'd5172,15'd5171,15'd5170,15'd5169,15'd5168,15'd5167,15'd5166,15'd5165,15'd5164,15'd5163,15'd5162,15'd5161,15'd5160,15'd5159,15'd5158,15'd5157,15'd5156,15'd5155,15'd5154,15'd5153,15'd5152,15'd5151,15'd5150,15'd5149,15'd5148,15'd5147,15'd5146,15'd5145,15'd5144,15'd5143,15'd5142,15'd5141,15'd5140,15'd5139,15'd5138,15'd5137,15'd5136,15'd5135,15'd5134,15'd5133,15'd5132,15'd5131,15'd5130,15'd5129,15'd5128,15'd5127,15'd5126,15'd5125,15'd5124,15'd5123,15'd5122,15'd5121,15'd5120,
15'd4879,15'd4878,15'd4877,15'd4876,15'd4875,15'd4874,15'd4873,15'd4872,15'd4871,15'd4870,15'd4869,15'd4868,15'd4867,15'd4866,15'd4865,15'd4864,15'd4863,15'd4862,15'd4861,15'd4860,15'd4859,15'd4858,15'd4857,15'd4856,15'd4855,15'd4854,15'd4853,15'd4852,15'd4851,15'd4850,15'd4849,15'd4848,15'd4847,15'd4846,15'd4845,15'd4844,15'd4843,15'd4842,15'd4841,15'd4840,15'd4839,15'd4838,15'd4837,15'd4836,15'd4835,15'd4834,15'd4833,15'd4832,15'd4831,15'd4830,15'd4829,15'd4828,15'd4827,15'd4826,15'd4825,15'd4824,15'd4823,15'd4822,15'd4821,15'd4820,15'd4819,15'd4818,15'd4817,15'd4816,15'd4815,15'd4814,15'd4813,15'd4812,15'd4811,15'd4810,15'd4809,15'd4808,15'd4807,15'd4806,15'd4805,15'd4804,15'd4803,15'd4802,15'd4801,15'd4800,
15'd4559,15'd4558,15'd4557,15'd4556,15'd4555,15'd4554,15'd4553,15'd4552,15'd4551,15'd4550,15'd4549,15'd4548,15'd4547,15'd4546,15'd4545,15'd4544,15'd4543,15'd4542,15'd4541,15'd4540,15'd4539,15'd4538,15'd4537,15'd4536,15'd4535,15'd4534,15'd4533,15'd4532,15'd4531,15'd4530,15'd4529,15'd4528,15'd4527,15'd4526,15'd4525,15'd4524,15'd4523,15'd4522,15'd4521,15'd4520,15'd4519,15'd4518,15'd4517,15'd4516,15'd4515,15'd4514,15'd4513,15'd4512,15'd4511,15'd4510,15'd4509,15'd4508,15'd4507,15'd4506,15'd4505,15'd4504,15'd4503,15'd4502,15'd4501,15'd4500,15'd4499,15'd4498,15'd4497,15'd4496,15'd4495,15'd4494,15'd4493,15'd4492,15'd4491,15'd4490,15'd4489,15'd4488,15'd4487,15'd4486,15'd4485,15'd4484,15'd4483,15'd4482,15'd4481,15'd4480,
15'd4239,15'd4238,15'd4237,15'd4236,15'd4235,15'd4234,15'd4233,15'd4232,15'd4231,15'd4230,15'd4229,15'd4228,15'd4227,15'd4226,15'd4225,15'd4224,15'd4223,15'd4222,15'd4221,15'd4220,15'd4219,15'd4218,15'd4217,15'd4216,15'd4215,15'd4214,15'd4213,15'd4212,15'd4211,15'd4210,15'd4209,15'd4208,15'd4207,15'd4206,15'd4205,15'd4204,15'd4203,15'd4202,15'd4201,15'd4200,15'd4199,15'd4198,15'd4197,15'd4196,15'd4195,15'd4194,15'd4193,15'd4192,15'd4191,15'd4190,15'd4189,15'd4188,15'd4187,15'd4186,15'd4185,15'd4184,15'd4183,15'd4182,15'd4181,15'd4180,15'd4179,15'd4178,15'd4177,15'd4176,15'd4175,15'd4174,15'd4173,15'd4172,15'd4171,15'd4170,15'd4169,15'd4168,15'd4167,15'd4166,15'd4165,15'd4164,15'd4163,15'd4162,15'd4161,15'd4160,
15'd3919,15'd3918,15'd3917,15'd3916,15'd3915,15'd3914,15'd3913,15'd3912,15'd3911,15'd3910,15'd3909,15'd3908,15'd3907,15'd3906,15'd3905,15'd3904,15'd3903,15'd3902,15'd3901,15'd3900,15'd3899,15'd3898,15'd3897,15'd3896,15'd3895,15'd3894,15'd3893,15'd3892,15'd3891,15'd3890,15'd3889,15'd3888,15'd3887,15'd3886,15'd3885,15'd3884,15'd3883,15'd3882,15'd3881,15'd3880,15'd3879,15'd3878,15'd3877,15'd3876,15'd3875,15'd3874,15'd3873,15'd3872,15'd3871,15'd3870,15'd3869,15'd3868,15'd3867,15'd3866,15'd3865,15'd3864,15'd3863,15'd3862,15'd3861,15'd3860,15'd3859,15'd3858,15'd3857,15'd3856,15'd3855,15'd3854,15'd3853,15'd3852,15'd3851,15'd3850,15'd3849,15'd3848,15'd3847,15'd3846,15'd3845,15'd3844,15'd3843,15'd3842,15'd3841,15'd3840,
15'd3599,15'd3598,15'd3597,15'd3596,15'd3595,15'd3594,15'd3593,15'd3592,15'd3591,15'd3590,15'd3589,15'd3588,15'd3587,15'd3586,15'd3585,15'd3584,15'd3583,15'd3582,15'd3581,15'd3580,15'd3579,15'd3578,15'd3577,15'd3576,15'd3575,15'd3574,15'd3573,15'd3572,15'd3571,15'd3570,15'd3569,15'd3568,15'd3567,15'd3566,15'd3565,15'd3564,15'd3563,15'd3562,15'd3561,15'd3560,15'd3559,15'd3558,15'd3557,15'd3556,15'd3555,15'd3554,15'd3553,15'd3552,15'd3551,15'd3550,15'd3549,15'd3548,15'd3547,15'd3546,15'd3545,15'd3544,15'd3543,15'd3542,15'd3541,15'd3540,15'd3539,15'd3538,15'd3537,15'd3536,15'd3535,15'd3534,15'd3533,15'd3532,15'd3531,15'd3530,15'd3529,15'd3528,15'd3527,15'd3526,15'd3525,15'd3524,15'd3523,15'd3522,15'd3521,15'd3520,
15'd3279,15'd3278,15'd3277,15'd3276,15'd3275,15'd3274,15'd3273,15'd3272,15'd3271,15'd3270,15'd3269,15'd3268,15'd3267,15'd3266,15'd3265,15'd3264,15'd3263,15'd3262,15'd3261,15'd3260,15'd3259,15'd3258,15'd3257,15'd3256,15'd3255,15'd3254,15'd3253,15'd3252,15'd3251,15'd3250,15'd3249,15'd3248,15'd3247,15'd3246,15'd3245,15'd3244,15'd3243,15'd3242,15'd3241,15'd3240,15'd3239,15'd3238,15'd3237,15'd3236,15'd3235,15'd3234,15'd3233,15'd3232,15'd3231,15'd3230,15'd3229,15'd3228,15'd3227,15'd3226,15'd3225,15'd3224,15'd3223,15'd3222,15'd3221,15'd3220,15'd3219,15'd3218,15'd3217,15'd3216,15'd3215,15'd3214,15'd3213,15'd3212,15'd3211,15'd3210,15'd3209,15'd3208,15'd3207,15'd3206,15'd3205,15'd3204,15'd3203,15'd3202,15'd3201,15'd3200,
15'd2959,15'd2958,15'd2957,15'd2956,15'd2955,15'd2954,15'd2953,15'd2952,15'd2951,15'd2950,15'd2949,15'd2948,15'd2947,15'd2946,15'd2945,15'd2944,15'd2943,15'd2942,15'd2941,15'd2940,15'd2939,15'd2938,15'd2937,15'd2936,15'd2935,15'd2934,15'd2933,15'd2932,15'd2931,15'd2930,15'd2929,15'd2928,15'd2927,15'd2926,15'd2925,15'd2924,15'd2923,15'd2922,15'd2921,15'd2920,15'd2919,15'd2918,15'd2917,15'd2916,15'd2915,15'd2914,15'd2913,15'd2912,15'd2911,15'd2910,15'd2909,15'd2908,15'd2907,15'd2906,15'd2905,15'd2904,15'd2903,15'd2902,15'd2901,15'd2900,15'd2899,15'd2898,15'd2897,15'd2896,15'd2895,15'd2894,15'd2893,15'd2892,15'd2891,15'd2890,15'd2889,15'd2888,15'd2887,15'd2886,15'd2885,15'd2884,15'd2883,15'd2882,15'd2881,15'd2880,
15'd2639,15'd2638,15'd2637,15'd2636,15'd2635,15'd2634,15'd2633,15'd2632,15'd2631,15'd2630,15'd2629,15'd2628,15'd2627,15'd2626,15'd2625,15'd2624,15'd2623,15'd2622,15'd2621,15'd2620,15'd2619,15'd2618,15'd2617,15'd2616,15'd2615,15'd2614,15'd2613,15'd2612,15'd2611,15'd2610,15'd2609,15'd2608,15'd2607,15'd2606,15'd2605,15'd2604,15'd2603,15'd2602,15'd2601,15'd2600,15'd2599,15'd2598,15'd2597,15'd2596,15'd2595,15'd2594,15'd2593,15'd2592,15'd2591,15'd2590,15'd2589,15'd2588,15'd2587,15'd2586,15'd2585,15'd2584,15'd2583,15'd2582,15'd2581,15'd2580,15'd2579,15'd2578,15'd2577,15'd2576,15'd2575,15'd2574,15'd2573,15'd2572,15'd2571,15'd2570,15'd2569,15'd2568,15'd2567,15'd2566,15'd2565,15'd2564,15'd2563,15'd2562,15'd2561,15'd2560,
15'd2319,15'd2318,15'd2317,15'd2316,15'd2315,15'd2314,15'd2313,15'd2312,15'd2311,15'd2310,15'd2309,15'd2308,15'd2307,15'd2306,15'd2305,15'd2304,15'd2303,15'd2302,15'd2301,15'd2300,15'd2299,15'd2298,15'd2297,15'd2296,15'd2295,15'd2294,15'd2293,15'd2292,15'd2291,15'd2290,15'd2289,15'd2288,15'd2287,15'd2286,15'd2285,15'd2284,15'd2283,15'd2282,15'd2281,15'd2280,15'd2279,15'd2278,15'd2277,15'd2276,15'd2275,15'd2274,15'd2273,15'd2272,15'd2271,15'd2270,15'd2269,15'd2268,15'd2267,15'd2266,15'd2265,15'd2264,15'd2263,15'd2262,15'd2261,15'd2260,15'd2259,15'd2258,15'd2257,15'd2256,15'd2255,15'd2254,15'd2253,15'd2252,15'd2251,15'd2250,15'd2249,15'd2248,15'd2247,15'd2246,15'd2245,15'd2244,15'd2243,15'd2242,15'd2241,15'd2240,
15'd1999,15'd1998,15'd1997,15'd1996,15'd1995,15'd1994,15'd1993,15'd1992,15'd1991,15'd1990,15'd1989,15'd1988,15'd1987,15'd1986,15'd1985,15'd1984,15'd1983,15'd1982,15'd1981,15'd1980,15'd1979,15'd1978,15'd1977,15'd1976,15'd1975,15'd1974,15'd1973,15'd1972,15'd1971,15'd1970,15'd1969,15'd1968,15'd1967,15'd1966,15'd1965,15'd1964,15'd1963,15'd1962,15'd1961,15'd1960,15'd1959,15'd1958,15'd1957,15'd1956,15'd1955,15'd1954,15'd1953,15'd1952,15'd1951,15'd1950,15'd1949,15'd1948,15'd1947,15'd1946,15'd1945,15'd1944,15'd1943,15'd1942,15'd1941,15'd1940,15'd1939,15'd1938,15'd1937,15'd1936,15'd1935,15'd1934,15'd1933,15'd1932,15'd1931,15'd1930,15'd1929,15'd1928,15'd1927,15'd1926,15'd1925,15'd1924,15'd1923,15'd1922,15'd1921,15'd1920,
15'd1679,15'd1678,15'd1677,15'd1676,15'd1675,15'd1674,15'd1673,15'd1672,15'd1671,15'd1670,15'd1669,15'd1668,15'd1667,15'd1666,15'd1665,15'd1664,15'd1663,15'd1662,15'd1661,15'd1660,15'd1659,15'd1658,15'd1657,15'd1656,15'd1655,15'd1654,15'd1653,15'd1652,15'd1651,15'd1650,15'd1649,15'd1648,15'd1647,15'd1646,15'd1645,15'd1644,15'd1643,15'd1642,15'd1641,15'd1640,15'd1639,15'd1638,15'd1637,15'd1636,15'd1635,15'd1634,15'd1633,15'd1632,15'd1631,15'd1630,15'd1629,15'd1628,15'd1627,15'd1626,15'd1625,15'd1624,15'd1623,15'd1622,15'd1621,15'd1620,15'd1619,15'd1618,15'd1617,15'd1616,15'd1615,15'd1614,15'd1613,15'd1612,15'd1611,15'd1610,15'd1609,15'd1608,15'd1607,15'd1606,15'd1605,15'd1604,15'd1603,15'd1602,15'd1601,15'd1600,
15'd1359,15'd1358,15'd1357,15'd1356,15'd1355,15'd1354,15'd1353,15'd1352,15'd1351,15'd1350,15'd1349,15'd1348,15'd1347,15'd1346,15'd1345,15'd1344,15'd1343,15'd1342,15'd1341,15'd1340,15'd1339,15'd1338,15'd1337,15'd1336,15'd1335,15'd1334,15'd1333,15'd1332,15'd1331,15'd1330,15'd1329,15'd1328,15'd1327,15'd1326,15'd1325,15'd1324,15'd1323,15'd1322,15'd1321,15'd1320,15'd1319,15'd1318,15'd1317,15'd1316,15'd1315,15'd1314,15'd1313,15'd1312,15'd1311,15'd1310,15'd1309,15'd1308,15'd1307,15'd1306,15'd1305,15'd1304,15'd1303,15'd1302,15'd1301,15'd1300,15'd1299,15'd1298,15'd1297,15'd1296,15'd1295,15'd1294,15'd1293,15'd1292,15'd1291,15'd1290,15'd1289,15'd1288,15'd1287,15'd1286,15'd1285,15'd1284,15'd1283,15'd1282,15'd1281,15'd1280,
15'd1039,15'd1038,15'd1037,15'd1036,15'd1035,15'd1034,15'd1033,15'd1032,15'd1031,15'd1030,15'd1029,15'd1028,15'd1027,15'd1026,15'd1025,15'd1024,15'd1023,15'd1022,15'd1021,15'd1020,15'd1019,15'd1018,15'd1017,15'd1016,15'd1015,15'd1014,15'd1013,15'd1012,15'd1011,15'd1010,15'd1009,15'd1008,15'd1007,15'd1006,15'd1005,15'd1004,15'd1003,15'd1002,15'd1001,15'd1000,15'd999,15'd998,15'd997,15'd996,15'd995,15'd994,15'd993,15'd992,15'd991,15'd990,15'd989,15'd988,15'd987,15'd986,15'd985,15'd984,15'd983,15'd982,15'd981,15'd980,15'd979,15'd978,15'd977,15'd976,15'd975,15'd974,15'd973,15'd972,15'd971,15'd970,15'd969,15'd968,15'd967,15'd966,15'd965,15'd964,15'd963,15'd962,15'd961,15'd960,
15'd719,15'd718,15'd717,15'd716,15'd715,15'd714,15'd713,15'd712,15'd711,15'd710,15'd709,15'd708,15'd707,15'd706,15'd705,15'd704,15'd703,15'd702,15'd701,15'd700,15'd699,15'd698,15'd697,15'd696,15'd695,15'd694,15'd693,15'd692,15'd691,15'd690,15'd689,15'd688,15'd687,15'd686,15'd685,15'd684,15'd683,15'd682,15'd681,15'd680,15'd679,15'd678,15'd677,15'd676,15'd675,15'd674,15'd673,15'd672,15'd671,15'd670,15'd669,15'd668,15'd667,15'd666,15'd665,15'd664,15'd663,15'd662,15'd661,15'd660,15'd659,15'd658,15'd657,15'd656,15'd655,15'd654,15'd653,15'd652,15'd651,15'd650,15'd649,15'd648,15'd647,15'd646,15'd645,15'd644,15'd643,15'd642,15'd641,15'd640,
15'd399,15'd398,15'd397,15'd396,15'd395,15'd394,15'd393,15'd392,15'd391,15'd390,15'd389,15'd388,15'd387,15'd386,15'd385,15'd384,15'd383,15'd382,15'd381,15'd380,15'd379,15'd378,15'd377,15'd376,15'd375,15'd374,15'd373,15'd372,15'd371,15'd370,15'd369,15'd368,15'd367,15'd366,15'd365,15'd364,15'd363,15'd362,15'd361,15'd360,15'd359,15'd358,15'd357,15'd356,15'd355,15'd354,15'd353,15'd352,15'd351,15'd350,15'd349,15'd348,15'd347,15'd346,15'd345,15'd344,15'd343,15'd342,15'd341,15'd340,15'd339,15'd338,15'd337,15'd336,15'd335,15'd334,15'd333,15'd332,15'd331,15'd330,15'd329,15'd328,15'd327,15'd326,15'd325,15'd324,15'd323,15'd322,15'd321,15'd320,
15'd79,15'd78,15'd77,15'd76,15'd75,15'd74,15'd73,15'd72,15'd71,15'd70,15'd69,15'd68,15'd67,15'd66,15'd65,15'd64,15'd63,15'd62,15'd61,15'd60,15'd59,15'd58,15'd57,15'd56,15'd55,15'd54,15'd53,15'd52,15'd51,15'd50,15'd49,15'd48,15'd47,15'd46,15'd45,15'd44,15'd43,15'd42,15'd41,15'd40,15'd39,15'd38,15'd37,15'd36,15'd35,15'd34,15'd33,15'd32,15'd31,15'd30,15'd29,15'd28,15'd27,15'd26,15'd25,15'd24,15'd23,15'd22,15'd21,15'd20,15'd19,15'd18,15'd17,15'd16,15'd15,15'd14,15'd13,15'd12,15'd11,15'd10,15'd9,15'd8,15'd7,15'd6,15'd5,15'd4,15'd3,15'd2,15'd1,15'd0};
parameter [14:0] state_3 [0:6399] = {
15'd79,15'd399,15'd719,15'd1039,15'd1359,15'd1679,15'd1999,15'd2319,15'd2639,15'd2959,15'd3279,15'd3599,15'd3919,15'd4239,15'd4559,15'd4879,15'd5199,15'd5519,15'd5839,15'd6159,15'd6479,15'd6799,15'd7119,15'd7439,15'd7759,15'd8079,15'd8399,15'd8719,15'd9039,15'd9359,15'd9679,15'd9999,15'd10319,15'd10639,15'd10959,15'd11279,15'd11599,15'd11919,15'd12239,15'd12559,15'd12879,15'd13199,15'd13519,15'd13839,15'd14159,15'd14479,15'd14799,15'd15119,15'd15439,15'd15759,15'd16079,15'd16399,15'd16719,15'd17039,15'd17359,15'd17679,15'd17999,15'd18319,15'd18639,15'd18959,15'd19279,15'd19599,15'd19919,15'd20239,15'd20559,15'd20879,15'd21199,15'd21519,15'd21839,15'd22159,15'd22479,15'd22799,15'd23119,15'd23439,15'd23759,15'd24079,15'd24399,15'd24719,15'd25039,15'd25359,
15'd78,15'd398,15'd718,15'd1038,15'd1358,15'd1678,15'd1998,15'd2318,15'd2638,15'd2958,15'd3278,15'd3598,15'd3918,15'd4238,15'd4558,15'd4878,15'd5198,15'd5518,15'd5838,15'd6158,15'd6478,15'd6798,15'd7118,15'd7438,15'd7758,15'd8078,15'd8398,15'd8718,15'd9038,15'd9358,15'd9678,15'd9998,15'd10318,15'd10638,15'd10958,15'd11278,15'd11598,15'd11918,15'd12238,15'd12558,15'd12878,15'd13198,15'd13518,15'd13838,15'd14158,15'd14478,15'd14798,15'd15118,15'd15438,15'd15758,15'd16078,15'd16398,15'd16718,15'd17038,15'd17358,15'd17678,15'd17998,15'd18318,15'd18638,15'd18958,15'd19278,15'd19598,15'd19918,15'd20238,15'd20558,15'd20878,15'd21198,15'd21518,15'd21838,15'd22158,15'd22478,15'd22798,15'd23118,15'd23438,15'd23758,15'd24078,15'd24398,15'd24718,15'd25038,15'd25358,
15'd77,15'd397,15'd717,15'd1037,15'd1357,15'd1677,15'd1997,15'd2317,15'd2637,15'd2957,15'd3277,15'd3597,15'd3917,15'd4237,15'd4557,15'd4877,15'd5197,15'd5517,15'd5837,15'd6157,15'd6477,15'd6797,15'd7117,15'd7437,15'd7757,15'd8077,15'd8397,15'd8717,15'd9037,15'd9357,15'd9677,15'd9997,15'd10317,15'd10637,15'd10957,15'd11277,15'd11597,15'd11917,15'd12237,15'd12557,15'd12877,15'd13197,15'd13517,15'd13837,15'd14157,15'd14477,15'd14797,15'd15117,15'd15437,15'd15757,15'd16077,15'd16397,15'd16717,15'd17037,15'd17357,15'd17677,15'd17997,15'd18317,15'd18637,15'd18957,15'd19277,15'd19597,15'd19917,15'd20237,15'd20557,15'd20877,15'd21197,15'd21517,15'd21837,15'd22157,15'd22477,15'd22797,15'd23117,15'd23437,15'd23757,15'd24077,15'd24397,15'd24717,15'd25037,15'd25357,
15'd76,15'd396,15'd716,15'd1036,15'd1356,15'd1676,15'd1996,15'd2316,15'd2636,15'd2956,15'd3276,15'd3596,15'd3916,15'd4236,15'd4556,15'd4876,15'd5196,15'd5516,15'd5836,15'd6156,15'd6476,15'd6796,15'd7116,15'd7436,15'd7756,15'd8076,15'd8396,15'd8716,15'd9036,15'd9356,15'd9676,15'd9996,15'd10316,15'd10636,15'd10956,15'd11276,15'd11596,15'd11916,15'd12236,15'd12556,15'd12876,15'd13196,15'd13516,15'd13836,15'd14156,15'd14476,15'd14796,15'd15116,15'd15436,15'd15756,15'd16076,15'd16396,15'd16716,15'd17036,15'd17356,15'd17676,15'd17996,15'd18316,15'd18636,15'd18956,15'd19276,15'd19596,15'd19916,15'd20236,15'd20556,15'd20876,15'd21196,15'd21516,15'd21836,15'd22156,15'd22476,15'd22796,15'd23116,15'd23436,15'd23756,15'd24076,15'd24396,15'd24716,15'd25036,15'd25356,
15'd75,15'd395,15'd715,15'd1035,15'd1355,15'd1675,15'd1995,15'd2315,15'd2635,15'd2955,15'd3275,15'd3595,15'd3915,15'd4235,15'd4555,15'd4875,15'd5195,15'd5515,15'd5835,15'd6155,15'd6475,15'd6795,15'd7115,15'd7435,15'd7755,15'd8075,15'd8395,15'd8715,15'd9035,15'd9355,15'd9675,15'd9995,15'd10315,15'd10635,15'd10955,15'd11275,15'd11595,15'd11915,15'd12235,15'd12555,15'd12875,15'd13195,15'd13515,15'd13835,15'd14155,15'd14475,15'd14795,15'd15115,15'd15435,15'd15755,15'd16075,15'd16395,15'd16715,15'd17035,15'd17355,15'd17675,15'd17995,15'd18315,15'd18635,15'd18955,15'd19275,15'd19595,15'd19915,15'd20235,15'd20555,15'd20875,15'd21195,15'd21515,15'd21835,15'd22155,15'd22475,15'd22795,15'd23115,15'd23435,15'd23755,15'd24075,15'd24395,15'd24715,15'd25035,15'd25355,
15'd74,15'd394,15'd714,15'd1034,15'd1354,15'd1674,15'd1994,15'd2314,15'd2634,15'd2954,15'd3274,15'd3594,15'd3914,15'd4234,15'd4554,15'd4874,15'd5194,15'd5514,15'd5834,15'd6154,15'd6474,15'd6794,15'd7114,15'd7434,15'd7754,15'd8074,15'd8394,15'd8714,15'd9034,15'd9354,15'd9674,15'd9994,15'd10314,15'd10634,15'd10954,15'd11274,15'd11594,15'd11914,15'd12234,15'd12554,15'd12874,15'd13194,15'd13514,15'd13834,15'd14154,15'd14474,15'd14794,15'd15114,15'd15434,15'd15754,15'd16074,15'd16394,15'd16714,15'd17034,15'd17354,15'd17674,15'd17994,15'd18314,15'd18634,15'd18954,15'd19274,15'd19594,15'd19914,15'd20234,15'd20554,15'd20874,15'd21194,15'd21514,15'd21834,15'd22154,15'd22474,15'd22794,15'd23114,15'd23434,15'd23754,15'd24074,15'd24394,15'd24714,15'd25034,15'd25354,
15'd73,15'd393,15'd713,15'd1033,15'd1353,15'd1673,15'd1993,15'd2313,15'd2633,15'd2953,15'd3273,15'd3593,15'd3913,15'd4233,15'd4553,15'd4873,15'd5193,15'd5513,15'd5833,15'd6153,15'd6473,15'd6793,15'd7113,15'd7433,15'd7753,15'd8073,15'd8393,15'd8713,15'd9033,15'd9353,15'd9673,15'd9993,15'd10313,15'd10633,15'd10953,15'd11273,15'd11593,15'd11913,15'd12233,15'd12553,15'd12873,15'd13193,15'd13513,15'd13833,15'd14153,15'd14473,15'd14793,15'd15113,15'd15433,15'd15753,15'd16073,15'd16393,15'd16713,15'd17033,15'd17353,15'd17673,15'd17993,15'd18313,15'd18633,15'd18953,15'd19273,15'd19593,15'd19913,15'd20233,15'd20553,15'd20873,15'd21193,15'd21513,15'd21833,15'd22153,15'd22473,15'd22793,15'd23113,15'd23433,15'd23753,15'd24073,15'd24393,15'd24713,15'd25033,15'd25353,
15'd72,15'd392,15'd712,15'd1032,15'd1352,15'd1672,15'd1992,15'd2312,15'd2632,15'd2952,15'd3272,15'd3592,15'd3912,15'd4232,15'd4552,15'd4872,15'd5192,15'd5512,15'd5832,15'd6152,15'd6472,15'd6792,15'd7112,15'd7432,15'd7752,15'd8072,15'd8392,15'd8712,15'd9032,15'd9352,15'd9672,15'd9992,15'd10312,15'd10632,15'd10952,15'd11272,15'd11592,15'd11912,15'd12232,15'd12552,15'd12872,15'd13192,15'd13512,15'd13832,15'd14152,15'd14472,15'd14792,15'd15112,15'd15432,15'd15752,15'd16072,15'd16392,15'd16712,15'd17032,15'd17352,15'd17672,15'd17992,15'd18312,15'd18632,15'd18952,15'd19272,15'd19592,15'd19912,15'd20232,15'd20552,15'd20872,15'd21192,15'd21512,15'd21832,15'd22152,15'd22472,15'd22792,15'd23112,15'd23432,15'd23752,15'd24072,15'd24392,15'd24712,15'd25032,15'd25352,
15'd71,15'd391,15'd711,15'd1031,15'd1351,15'd1671,15'd1991,15'd2311,15'd2631,15'd2951,15'd3271,15'd3591,15'd3911,15'd4231,15'd4551,15'd4871,15'd5191,15'd5511,15'd5831,15'd6151,15'd6471,15'd6791,15'd7111,15'd7431,15'd7751,15'd8071,15'd8391,15'd8711,15'd9031,15'd9351,15'd9671,15'd9991,15'd10311,15'd10631,15'd10951,15'd11271,15'd11591,15'd11911,15'd12231,15'd12551,15'd12871,15'd13191,15'd13511,15'd13831,15'd14151,15'd14471,15'd14791,15'd15111,15'd15431,15'd15751,15'd16071,15'd16391,15'd16711,15'd17031,15'd17351,15'd17671,15'd17991,15'd18311,15'd18631,15'd18951,15'd19271,15'd19591,15'd19911,15'd20231,15'd20551,15'd20871,15'd21191,15'd21511,15'd21831,15'd22151,15'd22471,15'd22791,15'd23111,15'd23431,15'd23751,15'd24071,15'd24391,15'd24711,15'd25031,15'd25351,
15'd70,15'd390,15'd710,15'd1030,15'd1350,15'd1670,15'd1990,15'd2310,15'd2630,15'd2950,15'd3270,15'd3590,15'd3910,15'd4230,15'd4550,15'd4870,15'd5190,15'd5510,15'd5830,15'd6150,15'd6470,15'd6790,15'd7110,15'd7430,15'd7750,15'd8070,15'd8390,15'd8710,15'd9030,15'd9350,15'd9670,15'd9990,15'd10310,15'd10630,15'd10950,15'd11270,15'd11590,15'd11910,15'd12230,15'd12550,15'd12870,15'd13190,15'd13510,15'd13830,15'd14150,15'd14470,15'd14790,15'd15110,15'd15430,15'd15750,15'd16070,15'd16390,15'd16710,15'd17030,15'd17350,15'd17670,15'd17990,15'd18310,15'd18630,15'd18950,15'd19270,15'd19590,15'd19910,15'd20230,15'd20550,15'd20870,15'd21190,15'd21510,15'd21830,15'd22150,15'd22470,15'd22790,15'd23110,15'd23430,15'd23750,15'd24070,15'd24390,15'd24710,15'd25030,15'd25350,
15'd69,15'd389,15'd709,15'd1029,15'd1349,15'd1669,15'd1989,15'd2309,15'd2629,15'd2949,15'd3269,15'd3589,15'd3909,15'd4229,15'd4549,15'd4869,15'd5189,15'd5509,15'd5829,15'd6149,15'd6469,15'd6789,15'd7109,15'd7429,15'd7749,15'd8069,15'd8389,15'd8709,15'd9029,15'd9349,15'd9669,15'd9989,15'd10309,15'd10629,15'd10949,15'd11269,15'd11589,15'd11909,15'd12229,15'd12549,15'd12869,15'd13189,15'd13509,15'd13829,15'd14149,15'd14469,15'd14789,15'd15109,15'd15429,15'd15749,15'd16069,15'd16389,15'd16709,15'd17029,15'd17349,15'd17669,15'd17989,15'd18309,15'd18629,15'd18949,15'd19269,15'd19589,15'd19909,15'd20229,15'd20549,15'd20869,15'd21189,15'd21509,15'd21829,15'd22149,15'd22469,15'd22789,15'd23109,15'd23429,15'd23749,15'd24069,15'd24389,15'd24709,15'd25029,15'd25349,
15'd68,15'd388,15'd708,15'd1028,15'd1348,15'd1668,15'd1988,15'd2308,15'd2628,15'd2948,15'd3268,15'd3588,15'd3908,15'd4228,15'd4548,15'd4868,15'd5188,15'd5508,15'd5828,15'd6148,15'd6468,15'd6788,15'd7108,15'd7428,15'd7748,15'd8068,15'd8388,15'd8708,15'd9028,15'd9348,15'd9668,15'd9988,15'd10308,15'd10628,15'd10948,15'd11268,15'd11588,15'd11908,15'd12228,15'd12548,15'd12868,15'd13188,15'd13508,15'd13828,15'd14148,15'd14468,15'd14788,15'd15108,15'd15428,15'd15748,15'd16068,15'd16388,15'd16708,15'd17028,15'd17348,15'd17668,15'd17988,15'd18308,15'd18628,15'd18948,15'd19268,15'd19588,15'd19908,15'd20228,15'd20548,15'd20868,15'd21188,15'd21508,15'd21828,15'd22148,15'd22468,15'd22788,15'd23108,15'd23428,15'd23748,15'd24068,15'd24388,15'd24708,15'd25028,15'd25348,
15'd67,15'd387,15'd707,15'd1027,15'd1347,15'd1667,15'd1987,15'd2307,15'd2627,15'd2947,15'd3267,15'd3587,15'd3907,15'd4227,15'd4547,15'd4867,15'd5187,15'd5507,15'd5827,15'd6147,15'd6467,15'd6787,15'd7107,15'd7427,15'd7747,15'd8067,15'd8387,15'd8707,15'd9027,15'd9347,15'd9667,15'd9987,15'd10307,15'd10627,15'd10947,15'd11267,15'd11587,15'd11907,15'd12227,15'd12547,15'd12867,15'd13187,15'd13507,15'd13827,15'd14147,15'd14467,15'd14787,15'd15107,15'd15427,15'd15747,15'd16067,15'd16387,15'd16707,15'd17027,15'd17347,15'd17667,15'd17987,15'd18307,15'd18627,15'd18947,15'd19267,15'd19587,15'd19907,15'd20227,15'd20547,15'd20867,15'd21187,15'd21507,15'd21827,15'd22147,15'd22467,15'd22787,15'd23107,15'd23427,15'd23747,15'd24067,15'd24387,15'd24707,15'd25027,15'd25347,
15'd66,15'd386,15'd706,15'd1026,15'd1346,15'd1666,15'd1986,15'd2306,15'd2626,15'd2946,15'd3266,15'd3586,15'd3906,15'd4226,15'd4546,15'd4866,15'd5186,15'd5506,15'd5826,15'd6146,15'd6466,15'd6786,15'd7106,15'd7426,15'd7746,15'd8066,15'd8386,15'd8706,15'd9026,15'd9346,15'd9666,15'd9986,15'd10306,15'd10626,15'd10946,15'd11266,15'd11586,15'd11906,15'd12226,15'd12546,15'd12866,15'd13186,15'd13506,15'd13826,15'd14146,15'd14466,15'd14786,15'd15106,15'd15426,15'd15746,15'd16066,15'd16386,15'd16706,15'd17026,15'd17346,15'd17666,15'd17986,15'd18306,15'd18626,15'd18946,15'd19266,15'd19586,15'd19906,15'd20226,15'd20546,15'd20866,15'd21186,15'd21506,15'd21826,15'd22146,15'd22466,15'd22786,15'd23106,15'd23426,15'd23746,15'd24066,15'd24386,15'd24706,15'd25026,15'd25346,
15'd65,15'd385,15'd705,15'd1025,15'd1345,15'd1665,15'd1985,15'd2305,15'd2625,15'd2945,15'd3265,15'd3585,15'd3905,15'd4225,15'd4545,15'd4865,15'd5185,15'd5505,15'd5825,15'd6145,15'd6465,15'd6785,15'd7105,15'd7425,15'd7745,15'd8065,15'd8385,15'd8705,15'd9025,15'd9345,15'd9665,15'd9985,15'd10305,15'd10625,15'd10945,15'd11265,15'd11585,15'd11905,15'd12225,15'd12545,15'd12865,15'd13185,15'd13505,15'd13825,15'd14145,15'd14465,15'd14785,15'd15105,15'd15425,15'd15745,15'd16065,15'd16385,15'd16705,15'd17025,15'd17345,15'd17665,15'd17985,15'd18305,15'd18625,15'd18945,15'd19265,15'd19585,15'd19905,15'd20225,15'd20545,15'd20865,15'd21185,15'd21505,15'd21825,15'd22145,15'd22465,15'd22785,15'd23105,15'd23425,15'd23745,15'd24065,15'd24385,15'd24705,15'd25025,15'd25345,
15'd64,15'd384,15'd704,15'd1024,15'd1344,15'd1664,15'd1984,15'd2304,15'd2624,15'd2944,15'd3264,15'd3584,15'd3904,15'd4224,15'd4544,15'd4864,15'd5184,15'd5504,15'd5824,15'd6144,15'd6464,15'd6784,15'd7104,15'd7424,15'd7744,15'd8064,15'd8384,15'd8704,15'd9024,15'd9344,15'd9664,15'd9984,15'd10304,15'd10624,15'd10944,15'd11264,15'd11584,15'd11904,15'd12224,15'd12544,15'd12864,15'd13184,15'd13504,15'd13824,15'd14144,15'd14464,15'd14784,15'd15104,15'd15424,15'd15744,15'd16064,15'd16384,15'd16704,15'd17024,15'd17344,15'd17664,15'd17984,15'd18304,15'd18624,15'd18944,15'd19264,15'd19584,15'd19904,15'd20224,15'd20544,15'd20864,15'd21184,15'd21504,15'd21824,15'd22144,15'd22464,15'd22784,15'd23104,15'd23424,15'd23744,15'd24064,15'd24384,15'd24704,15'd25024,15'd25344,
15'd63,15'd383,15'd703,15'd1023,15'd1343,15'd1663,15'd1983,15'd2303,15'd2623,15'd2943,15'd3263,15'd3583,15'd3903,15'd4223,15'd4543,15'd4863,15'd5183,15'd5503,15'd5823,15'd6143,15'd6463,15'd6783,15'd7103,15'd7423,15'd7743,15'd8063,15'd8383,15'd8703,15'd9023,15'd9343,15'd9663,15'd9983,15'd10303,15'd10623,15'd10943,15'd11263,15'd11583,15'd11903,15'd12223,15'd12543,15'd12863,15'd13183,15'd13503,15'd13823,15'd14143,15'd14463,15'd14783,15'd15103,15'd15423,15'd15743,15'd16063,15'd16383,15'd16703,15'd17023,15'd17343,15'd17663,15'd17983,15'd18303,15'd18623,15'd18943,15'd19263,15'd19583,15'd19903,15'd20223,15'd20543,15'd20863,15'd21183,15'd21503,15'd21823,15'd22143,15'd22463,15'd22783,15'd23103,15'd23423,15'd23743,15'd24063,15'd24383,15'd24703,15'd25023,15'd25343,
15'd62,15'd382,15'd702,15'd1022,15'd1342,15'd1662,15'd1982,15'd2302,15'd2622,15'd2942,15'd3262,15'd3582,15'd3902,15'd4222,15'd4542,15'd4862,15'd5182,15'd5502,15'd5822,15'd6142,15'd6462,15'd6782,15'd7102,15'd7422,15'd7742,15'd8062,15'd8382,15'd8702,15'd9022,15'd9342,15'd9662,15'd9982,15'd10302,15'd10622,15'd10942,15'd11262,15'd11582,15'd11902,15'd12222,15'd12542,15'd12862,15'd13182,15'd13502,15'd13822,15'd14142,15'd14462,15'd14782,15'd15102,15'd15422,15'd15742,15'd16062,15'd16382,15'd16702,15'd17022,15'd17342,15'd17662,15'd17982,15'd18302,15'd18622,15'd18942,15'd19262,15'd19582,15'd19902,15'd20222,15'd20542,15'd20862,15'd21182,15'd21502,15'd21822,15'd22142,15'd22462,15'd22782,15'd23102,15'd23422,15'd23742,15'd24062,15'd24382,15'd24702,15'd25022,15'd25342,
15'd61,15'd381,15'd701,15'd1021,15'd1341,15'd1661,15'd1981,15'd2301,15'd2621,15'd2941,15'd3261,15'd3581,15'd3901,15'd4221,15'd4541,15'd4861,15'd5181,15'd5501,15'd5821,15'd6141,15'd6461,15'd6781,15'd7101,15'd7421,15'd7741,15'd8061,15'd8381,15'd8701,15'd9021,15'd9341,15'd9661,15'd9981,15'd10301,15'd10621,15'd10941,15'd11261,15'd11581,15'd11901,15'd12221,15'd12541,15'd12861,15'd13181,15'd13501,15'd13821,15'd14141,15'd14461,15'd14781,15'd15101,15'd15421,15'd15741,15'd16061,15'd16381,15'd16701,15'd17021,15'd17341,15'd17661,15'd17981,15'd18301,15'd18621,15'd18941,15'd19261,15'd19581,15'd19901,15'd20221,15'd20541,15'd20861,15'd21181,15'd21501,15'd21821,15'd22141,15'd22461,15'd22781,15'd23101,15'd23421,15'd23741,15'd24061,15'd24381,15'd24701,15'd25021,15'd25341,
15'd60,15'd380,15'd700,15'd1020,15'd1340,15'd1660,15'd1980,15'd2300,15'd2620,15'd2940,15'd3260,15'd3580,15'd3900,15'd4220,15'd4540,15'd4860,15'd5180,15'd5500,15'd5820,15'd6140,15'd6460,15'd6780,15'd7100,15'd7420,15'd7740,15'd8060,15'd8380,15'd8700,15'd9020,15'd9340,15'd9660,15'd9980,15'd10300,15'd10620,15'd10940,15'd11260,15'd11580,15'd11900,15'd12220,15'd12540,15'd12860,15'd13180,15'd13500,15'd13820,15'd14140,15'd14460,15'd14780,15'd15100,15'd15420,15'd15740,15'd16060,15'd16380,15'd16700,15'd17020,15'd17340,15'd17660,15'd17980,15'd18300,15'd18620,15'd18940,15'd19260,15'd19580,15'd19900,15'd20220,15'd20540,15'd20860,15'd21180,15'd21500,15'd21820,15'd22140,15'd22460,15'd22780,15'd23100,15'd23420,15'd23740,15'd24060,15'd24380,15'd24700,15'd25020,15'd25340,
15'd59,15'd379,15'd699,15'd1019,15'd1339,15'd1659,15'd1979,15'd2299,15'd2619,15'd2939,15'd3259,15'd3579,15'd3899,15'd4219,15'd4539,15'd4859,15'd5179,15'd5499,15'd5819,15'd6139,15'd6459,15'd6779,15'd7099,15'd7419,15'd7739,15'd8059,15'd8379,15'd8699,15'd9019,15'd9339,15'd9659,15'd9979,15'd10299,15'd10619,15'd10939,15'd11259,15'd11579,15'd11899,15'd12219,15'd12539,15'd12859,15'd13179,15'd13499,15'd13819,15'd14139,15'd14459,15'd14779,15'd15099,15'd15419,15'd15739,15'd16059,15'd16379,15'd16699,15'd17019,15'd17339,15'd17659,15'd17979,15'd18299,15'd18619,15'd18939,15'd19259,15'd19579,15'd19899,15'd20219,15'd20539,15'd20859,15'd21179,15'd21499,15'd21819,15'd22139,15'd22459,15'd22779,15'd23099,15'd23419,15'd23739,15'd24059,15'd24379,15'd24699,15'd25019,15'd25339,
15'd58,15'd378,15'd698,15'd1018,15'd1338,15'd1658,15'd1978,15'd2298,15'd2618,15'd2938,15'd3258,15'd3578,15'd3898,15'd4218,15'd4538,15'd4858,15'd5178,15'd5498,15'd5818,15'd6138,15'd6458,15'd6778,15'd7098,15'd7418,15'd7738,15'd8058,15'd8378,15'd8698,15'd9018,15'd9338,15'd9658,15'd9978,15'd10298,15'd10618,15'd10938,15'd11258,15'd11578,15'd11898,15'd12218,15'd12538,15'd12858,15'd13178,15'd13498,15'd13818,15'd14138,15'd14458,15'd14778,15'd15098,15'd15418,15'd15738,15'd16058,15'd16378,15'd16698,15'd17018,15'd17338,15'd17658,15'd17978,15'd18298,15'd18618,15'd18938,15'd19258,15'd19578,15'd19898,15'd20218,15'd20538,15'd20858,15'd21178,15'd21498,15'd21818,15'd22138,15'd22458,15'd22778,15'd23098,15'd23418,15'd23738,15'd24058,15'd24378,15'd24698,15'd25018,15'd25338,
15'd57,15'd377,15'd697,15'd1017,15'd1337,15'd1657,15'd1977,15'd2297,15'd2617,15'd2937,15'd3257,15'd3577,15'd3897,15'd4217,15'd4537,15'd4857,15'd5177,15'd5497,15'd5817,15'd6137,15'd6457,15'd6777,15'd7097,15'd7417,15'd7737,15'd8057,15'd8377,15'd8697,15'd9017,15'd9337,15'd9657,15'd9977,15'd10297,15'd10617,15'd10937,15'd11257,15'd11577,15'd11897,15'd12217,15'd12537,15'd12857,15'd13177,15'd13497,15'd13817,15'd14137,15'd14457,15'd14777,15'd15097,15'd15417,15'd15737,15'd16057,15'd16377,15'd16697,15'd17017,15'd17337,15'd17657,15'd17977,15'd18297,15'd18617,15'd18937,15'd19257,15'd19577,15'd19897,15'd20217,15'd20537,15'd20857,15'd21177,15'd21497,15'd21817,15'd22137,15'd22457,15'd22777,15'd23097,15'd23417,15'd23737,15'd24057,15'd24377,15'd24697,15'd25017,15'd25337,
15'd56,15'd376,15'd696,15'd1016,15'd1336,15'd1656,15'd1976,15'd2296,15'd2616,15'd2936,15'd3256,15'd3576,15'd3896,15'd4216,15'd4536,15'd4856,15'd5176,15'd5496,15'd5816,15'd6136,15'd6456,15'd6776,15'd7096,15'd7416,15'd7736,15'd8056,15'd8376,15'd8696,15'd9016,15'd9336,15'd9656,15'd9976,15'd10296,15'd10616,15'd10936,15'd11256,15'd11576,15'd11896,15'd12216,15'd12536,15'd12856,15'd13176,15'd13496,15'd13816,15'd14136,15'd14456,15'd14776,15'd15096,15'd15416,15'd15736,15'd16056,15'd16376,15'd16696,15'd17016,15'd17336,15'd17656,15'd17976,15'd18296,15'd18616,15'd18936,15'd19256,15'd19576,15'd19896,15'd20216,15'd20536,15'd20856,15'd21176,15'd21496,15'd21816,15'd22136,15'd22456,15'd22776,15'd23096,15'd23416,15'd23736,15'd24056,15'd24376,15'd24696,15'd25016,15'd25336,
15'd55,15'd375,15'd695,15'd1015,15'd1335,15'd1655,15'd1975,15'd2295,15'd2615,15'd2935,15'd3255,15'd3575,15'd3895,15'd4215,15'd4535,15'd4855,15'd5175,15'd5495,15'd5815,15'd6135,15'd6455,15'd6775,15'd7095,15'd7415,15'd7735,15'd8055,15'd8375,15'd8695,15'd9015,15'd9335,15'd9655,15'd9975,15'd10295,15'd10615,15'd10935,15'd11255,15'd11575,15'd11895,15'd12215,15'd12535,15'd12855,15'd13175,15'd13495,15'd13815,15'd14135,15'd14455,15'd14775,15'd15095,15'd15415,15'd15735,15'd16055,15'd16375,15'd16695,15'd17015,15'd17335,15'd17655,15'd17975,15'd18295,15'd18615,15'd18935,15'd19255,15'd19575,15'd19895,15'd20215,15'd20535,15'd20855,15'd21175,15'd21495,15'd21815,15'd22135,15'd22455,15'd22775,15'd23095,15'd23415,15'd23735,15'd24055,15'd24375,15'd24695,15'd25015,15'd25335,
15'd54,15'd374,15'd694,15'd1014,15'd1334,15'd1654,15'd1974,15'd2294,15'd2614,15'd2934,15'd3254,15'd3574,15'd3894,15'd4214,15'd4534,15'd4854,15'd5174,15'd5494,15'd5814,15'd6134,15'd6454,15'd6774,15'd7094,15'd7414,15'd7734,15'd8054,15'd8374,15'd8694,15'd9014,15'd9334,15'd9654,15'd9974,15'd10294,15'd10614,15'd10934,15'd11254,15'd11574,15'd11894,15'd12214,15'd12534,15'd12854,15'd13174,15'd13494,15'd13814,15'd14134,15'd14454,15'd14774,15'd15094,15'd15414,15'd15734,15'd16054,15'd16374,15'd16694,15'd17014,15'd17334,15'd17654,15'd17974,15'd18294,15'd18614,15'd18934,15'd19254,15'd19574,15'd19894,15'd20214,15'd20534,15'd20854,15'd21174,15'd21494,15'd21814,15'd22134,15'd22454,15'd22774,15'd23094,15'd23414,15'd23734,15'd24054,15'd24374,15'd24694,15'd25014,15'd25334,
15'd53,15'd373,15'd693,15'd1013,15'd1333,15'd1653,15'd1973,15'd2293,15'd2613,15'd2933,15'd3253,15'd3573,15'd3893,15'd4213,15'd4533,15'd4853,15'd5173,15'd5493,15'd5813,15'd6133,15'd6453,15'd6773,15'd7093,15'd7413,15'd7733,15'd8053,15'd8373,15'd8693,15'd9013,15'd9333,15'd9653,15'd9973,15'd10293,15'd10613,15'd10933,15'd11253,15'd11573,15'd11893,15'd12213,15'd12533,15'd12853,15'd13173,15'd13493,15'd13813,15'd14133,15'd14453,15'd14773,15'd15093,15'd15413,15'd15733,15'd16053,15'd16373,15'd16693,15'd17013,15'd17333,15'd17653,15'd17973,15'd18293,15'd18613,15'd18933,15'd19253,15'd19573,15'd19893,15'd20213,15'd20533,15'd20853,15'd21173,15'd21493,15'd21813,15'd22133,15'd22453,15'd22773,15'd23093,15'd23413,15'd23733,15'd24053,15'd24373,15'd24693,15'd25013,15'd25333,
15'd52,15'd372,15'd692,15'd1012,15'd1332,15'd1652,15'd1972,15'd2292,15'd2612,15'd2932,15'd3252,15'd3572,15'd3892,15'd4212,15'd4532,15'd4852,15'd5172,15'd5492,15'd5812,15'd6132,15'd6452,15'd6772,15'd7092,15'd7412,15'd7732,15'd8052,15'd8372,15'd8692,15'd9012,15'd9332,15'd9652,15'd9972,15'd10292,15'd10612,15'd10932,15'd11252,15'd11572,15'd11892,15'd12212,15'd12532,15'd12852,15'd13172,15'd13492,15'd13812,15'd14132,15'd14452,15'd14772,15'd15092,15'd15412,15'd15732,15'd16052,15'd16372,15'd16692,15'd17012,15'd17332,15'd17652,15'd17972,15'd18292,15'd18612,15'd18932,15'd19252,15'd19572,15'd19892,15'd20212,15'd20532,15'd20852,15'd21172,15'd21492,15'd21812,15'd22132,15'd22452,15'd22772,15'd23092,15'd23412,15'd23732,15'd24052,15'd24372,15'd24692,15'd25012,15'd25332,
15'd51,15'd371,15'd691,15'd1011,15'd1331,15'd1651,15'd1971,15'd2291,15'd2611,15'd2931,15'd3251,15'd3571,15'd3891,15'd4211,15'd4531,15'd4851,15'd5171,15'd5491,15'd5811,15'd6131,15'd6451,15'd6771,15'd7091,15'd7411,15'd7731,15'd8051,15'd8371,15'd8691,15'd9011,15'd9331,15'd9651,15'd9971,15'd10291,15'd10611,15'd10931,15'd11251,15'd11571,15'd11891,15'd12211,15'd12531,15'd12851,15'd13171,15'd13491,15'd13811,15'd14131,15'd14451,15'd14771,15'd15091,15'd15411,15'd15731,15'd16051,15'd16371,15'd16691,15'd17011,15'd17331,15'd17651,15'd17971,15'd18291,15'd18611,15'd18931,15'd19251,15'd19571,15'd19891,15'd20211,15'd20531,15'd20851,15'd21171,15'd21491,15'd21811,15'd22131,15'd22451,15'd22771,15'd23091,15'd23411,15'd23731,15'd24051,15'd24371,15'd24691,15'd25011,15'd25331,
15'd50,15'd370,15'd690,15'd1010,15'd1330,15'd1650,15'd1970,15'd2290,15'd2610,15'd2930,15'd3250,15'd3570,15'd3890,15'd4210,15'd4530,15'd4850,15'd5170,15'd5490,15'd5810,15'd6130,15'd6450,15'd6770,15'd7090,15'd7410,15'd7730,15'd8050,15'd8370,15'd8690,15'd9010,15'd9330,15'd9650,15'd9970,15'd10290,15'd10610,15'd10930,15'd11250,15'd11570,15'd11890,15'd12210,15'd12530,15'd12850,15'd13170,15'd13490,15'd13810,15'd14130,15'd14450,15'd14770,15'd15090,15'd15410,15'd15730,15'd16050,15'd16370,15'd16690,15'd17010,15'd17330,15'd17650,15'd17970,15'd18290,15'd18610,15'd18930,15'd19250,15'd19570,15'd19890,15'd20210,15'd20530,15'd20850,15'd21170,15'd21490,15'd21810,15'd22130,15'd22450,15'd22770,15'd23090,15'd23410,15'd23730,15'd24050,15'd24370,15'd24690,15'd25010,15'd25330,
15'd49,15'd369,15'd689,15'd1009,15'd1329,15'd1649,15'd1969,15'd2289,15'd2609,15'd2929,15'd3249,15'd3569,15'd3889,15'd4209,15'd4529,15'd4849,15'd5169,15'd5489,15'd5809,15'd6129,15'd6449,15'd6769,15'd7089,15'd7409,15'd7729,15'd8049,15'd8369,15'd8689,15'd9009,15'd9329,15'd9649,15'd9969,15'd10289,15'd10609,15'd10929,15'd11249,15'd11569,15'd11889,15'd12209,15'd12529,15'd12849,15'd13169,15'd13489,15'd13809,15'd14129,15'd14449,15'd14769,15'd15089,15'd15409,15'd15729,15'd16049,15'd16369,15'd16689,15'd17009,15'd17329,15'd17649,15'd17969,15'd18289,15'd18609,15'd18929,15'd19249,15'd19569,15'd19889,15'd20209,15'd20529,15'd20849,15'd21169,15'd21489,15'd21809,15'd22129,15'd22449,15'd22769,15'd23089,15'd23409,15'd23729,15'd24049,15'd24369,15'd24689,15'd25009,15'd25329,
15'd48,15'd368,15'd688,15'd1008,15'd1328,15'd1648,15'd1968,15'd2288,15'd2608,15'd2928,15'd3248,15'd3568,15'd3888,15'd4208,15'd4528,15'd4848,15'd5168,15'd5488,15'd5808,15'd6128,15'd6448,15'd6768,15'd7088,15'd7408,15'd7728,15'd8048,15'd8368,15'd8688,15'd9008,15'd9328,15'd9648,15'd9968,15'd10288,15'd10608,15'd10928,15'd11248,15'd11568,15'd11888,15'd12208,15'd12528,15'd12848,15'd13168,15'd13488,15'd13808,15'd14128,15'd14448,15'd14768,15'd15088,15'd15408,15'd15728,15'd16048,15'd16368,15'd16688,15'd17008,15'd17328,15'd17648,15'd17968,15'd18288,15'd18608,15'd18928,15'd19248,15'd19568,15'd19888,15'd20208,15'd20528,15'd20848,15'd21168,15'd21488,15'd21808,15'd22128,15'd22448,15'd22768,15'd23088,15'd23408,15'd23728,15'd24048,15'd24368,15'd24688,15'd25008,15'd25328,
15'd47,15'd367,15'd687,15'd1007,15'd1327,15'd1647,15'd1967,15'd2287,15'd2607,15'd2927,15'd3247,15'd3567,15'd3887,15'd4207,15'd4527,15'd4847,15'd5167,15'd5487,15'd5807,15'd6127,15'd6447,15'd6767,15'd7087,15'd7407,15'd7727,15'd8047,15'd8367,15'd8687,15'd9007,15'd9327,15'd9647,15'd9967,15'd10287,15'd10607,15'd10927,15'd11247,15'd11567,15'd11887,15'd12207,15'd12527,15'd12847,15'd13167,15'd13487,15'd13807,15'd14127,15'd14447,15'd14767,15'd15087,15'd15407,15'd15727,15'd16047,15'd16367,15'd16687,15'd17007,15'd17327,15'd17647,15'd17967,15'd18287,15'd18607,15'd18927,15'd19247,15'd19567,15'd19887,15'd20207,15'd20527,15'd20847,15'd21167,15'd21487,15'd21807,15'd22127,15'd22447,15'd22767,15'd23087,15'd23407,15'd23727,15'd24047,15'd24367,15'd24687,15'd25007,15'd25327,
15'd46,15'd366,15'd686,15'd1006,15'd1326,15'd1646,15'd1966,15'd2286,15'd2606,15'd2926,15'd3246,15'd3566,15'd3886,15'd4206,15'd4526,15'd4846,15'd5166,15'd5486,15'd5806,15'd6126,15'd6446,15'd6766,15'd7086,15'd7406,15'd7726,15'd8046,15'd8366,15'd8686,15'd9006,15'd9326,15'd9646,15'd9966,15'd10286,15'd10606,15'd10926,15'd11246,15'd11566,15'd11886,15'd12206,15'd12526,15'd12846,15'd13166,15'd13486,15'd13806,15'd14126,15'd14446,15'd14766,15'd15086,15'd15406,15'd15726,15'd16046,15'd16366,15'd16686,15'd17006,15'd17326,15'd17646,15'd17966,15'd18286,15'd18606,15'd18926,15'd19246,15'd19566,15'd19886,15'd20206,15'd20526,15'd20846,15'd21166,15'd21486,15'd21806,15'd22126,15'd22446,15'd22766,15'd23086,15'd23406,15'd23726,15'd24046,15'd24366,15'd24686,15'd25006,15'd25326,
15'd45,15'd365,15'd685,15'd1005,15'd1325,15'd1645,15'd1965,15'd2285,15'd2605,15'd2925,15'd3245,15'd3565,15'd3885,15'd4205,15'd4525,15'd4845,15'd5165,15'd5485,15'd5805,15'd6125,15'd6445,15'd6765,15'd7085,15'd7405,15'd7725,15'd8045,15'd8365,15'd8685,15'd9005,15'd9325,15'd9645,15'd9965,15'd10285,15'd10605,15'd10925,15'd11245,15'd11565,15'd11885,15'd12205,15'd12525,15'd12845,15'd13165,15'd13485,15'd13805,15'd14125,15'd14445,15'd14765,15'd15085,15'd15405,15'd15725,15'd16045,15'd16365,15'd16685,15'd17005,15'd17325,15'd17645,15'd17965,15'd18285,15'd18605,15'd18925,15'd19245,15'd19565,15'd19885,15'd20205,15'd20525,15'd20845,15'd21165,15'd21485,15'd21805,15'd22125,15'd22445,15'd22765,15'd23085,15'd23405,15'd23725,15'd24045,15'd24365,15'd24685,15'd25005,15'd25325,
15'd44,15'd364,15'd684,15'd1004,15'd1324,15'd1644,15'd1964,15'd2284,15'd2604,15'd2924,15'd3244,15'd3564,15'd3884,15'd4204,15'd4524,15'd4844,15'd5164,15'd5484,15'd5804,15'd6124,15'd6444,15'd6764,15'd7084,15'd7404,15'd7724,15'd8044,15'd8364,15'd8684,15'd9004,15'd9324,15'd9644,15'd9964,15'd10284,15'd10604,15'd10924,15'd11244,15'd11564,15'd11884,15'd12204,15'd12524,15'd12844,15'd13164,15'd13484,15'd13804,15'd14124,15'd14444,15'd14764,15'd15084,15'd15404,15'd15724,15'd16044,15'd16364,15'd16684,15'd17004,15'd17324,15'd17644,15'd17964,15'd18284,15'd18604,15'd18924,15'd19244,15'd19564,15'd19884,15'd20204,15'd20524,15'd20844,15'd21164,15'd21484,15'd21804,15'd22124,15'd22444,15'd22764,15'd23084,15'd23404,15'd23724,15'd24044,15'd24364,15'd24684,15'd25004,15'd25324,
15'd43,15'd363,15'd683,15'd1003,15'd1323,15'd1643,15'd1963,15'd2283,15'd2603,15'd2923,15'd3243,15'd3563,15'd3883,15'd4203,15'd4523,15'd4843,15'd5163,15'd5483,15'd5803,15'd6123,15'd6443,15'd6763,15'd7083,15'd7403,15'd7723,15'd8043,15'd8363,15'd8683,15'd9003,15'd9323,15'd9643,15'd9963,15'd10283,15'd10603,15'd10923,15'd11243,15'd11563,15'd11883,15'd12203,15'd12523,15'd12843,15'd13163,15'd13483,15'd13803,15'd14123,15'd14443,15'd14763,15'd15083,15'd15403,15'd15723,15'd16043,15'd16363,15'd16683,15'd17003,15'd17323,15'd17643,15'd17963,15'd18283,15'd18603,15'd18923,15'd19243,15'd19563,15'd19883,15'd20203,15'd20523,15'd20843,15'd21163,15'd21483,15'd21803,15'd22123,15'd22443,15'd22763,15'd23083,15'd23403,15'd23723,15'd24043,15'd24363,15'd24683,15'd25003,15'd25323,
15'd42,15'd362,15'd682,15'd1002,15'd1322,15'd1642,15'd1962,15'd2282,15'd2602,15'd2922,15'd3242,15'd3562,15'd3882,15'd4202,15'd4522,15'd4842,15'd5162,15'd5482,15'd5802,15'd6122,15'd6442,15'd6762,15'd7082,15'd7402,15'd7722,15'd8042,15'd8362,15'd8682,15'd9002,15'd9322,15'd9642,15'd9962,15'd10282,15'd10602,15'd10922,15'd11242,15'd11562,15'd11882,15'd12202,15'd12522,15'd12842,15'd13162,15'd13482,15'd13802,15'd14122,15'd14442,15'd14762,15'd15082,15'd15402,15'd15722,15'd16042,15'd16362,15'd16682,15'd17002,15'd17322,15'd17642,15'd17962,15'd18282,15'd18602,15'd18922,15'd19242,15'd19562,15'd19882,15'd20202,15'd20522,15'd20842,15'd21162,15'd21482,15'd21802,15'd22122,15'd22442,15'd22762,15'd23082,15'd23402,15'd23722,15'd24042,15'd24362,15'd24682,15'd25002,15'd25322,
15'd41,15'd361,15'd681,15'd1001,15'd1321,15'd1641,15'd1961,15'd2281,15'd2601,15'd2921,15'd3241,15'd3561,15'd3881,15'd4201,15'd4521,15'd4841,15'd5161,15'd5481,15'd5801,15'd6121,15'd6441,15'd6761,15'd7081,15'd7401,15'd7721,15'd8041,15'd8361,15'd8681,15'd9001,15'd9321,15'd9641,15'd9961,15'd10281,15'd10601,15'd10921,15'd11241,15'd11561,15'd11881,15'd12201,15'd12521,15'd12841,15'd13161,15'd13481,15'd13801,15'd14121,15'd14441,15'd14761,15'd15081,15'd15401,15'd15721,15'd16041,15'd16361,15'd16681,15'd17001,15'd17321,15'd17641,15'd17961,15'd18281,15'd18601,15'd18921,15'd19241,15'd19561,15'd19881,15'd20201,15'd20521,15'd20841,15'd21161,15'd21481,15'd21801,15'd22121,15'd22441,15'd22761,15'd23081,15'd23401,15'd23721,15'd24041,15'd24361,15'd24681,15'd25001,15'd25321,
15'd40,15'd360,15'd680,15'd1000,15'd1320,15'd1640,15'd1960,15'd2280,15'd2600,15'd2920,15'd3240,15'd3560,15'd3880,15'd4200,15'd4520,15'd4840,15'd5160,15'd5480,15'd5800,15'd6120,15'd6440,15'd6760,15'd7080,15'd7400,15'd7720,15'd8040,15'd8360,15'd8680,15'd9000,15'd9320,15'd9640,15'd9960,15'd10280,15'd10600,15'd10920,15'd11240,15'd11560,15'd11880,15'd12200,15'd12520,15'd12840,15'd13160,15'd13480,15'd13800,15'd14120,15'd14440,15'd14760,15'd15080,15'd15400,15'd15720,15'd16040,15'd16360,15'd16680,15'd17000,15'd17320,15'd17640,15'd17960,15'd18280,15'd18600,15'd18920,15'd19240,15'd19560,15'd19880,15'd20200,15'd20520,15'd20840,15'd21160,15'd21480,15'd21800,15'd22120,15'd22440,15'd22760,15'd23080,15'd23400,15'd23720,15'd24040,15'd24360,15'd24680,15'd25000,15'd25320,
15'd39,15'd359,15'd679,15'd999,15'd1319,15'd1639,15'd1959,15'd2279,15'd2599,15'd2919,15'd3239,15'd3559,15'd3879,15'd4199,15'd4519,15'd4839,15'd5159,15'd5479,15'd5799,15'd6119,15'd6439,15'd6759,15'd7079,15'd7399,15'd7719,15'd8039,15'd8359,15'd8679,15'd8999,15'd9319,15'd9639,15'd9959,15'd10279,15'd10599,15'd10919,15'd11239,15'd11559,15'd11879,15'd12199,15'd12519,15'd12839,15'd13159,15'd13479,15'd13799,15'd14119,15'd14439,15'd14759,15'd15079,15'd15399,15'd15719,15'd16039,15'd16359,15'd16679,15'd16999,15'd17319,15'd17639,15'd17959,15'd18279,15'd18599,15'd18919,15'd19239,15'd19559,15'd19879,15'd20199,15'd20519,15'd20839,15'd21159,15'd21479,15'd21799,15'd22119,15'd22439,15'd22759,15'd23079,15'd23399,15'd23719,15'd24039,15'd24359,15'd24679,15'd24999,15'd25319,
15'd38,15'd358,15'd678,15'd998,15'd1318,15'd1638,15'd1958,15'd2278,15'd2598,15'd2918,15'd3238,15'd3558,15'd3878,15'd4198,15'd4518,15'd4838,15'd5158,15'd5478,15'd5798,15'd6118,15'd6438,15'd6758,15'd7078,15'd7398,15'd7718,15'd8038,15'd8358,15'd8678,15'd8998,15'd9318,15'd9638,15'd9958,15'd10278,15'd10598,15'd10918,15'd11238,15'd11558,15'd11878,15'd12198,15'd12518,15'd12838,15'd13158,15'd13478,15'd13798,15'd14118,15'd14438,15'd14758,15'd15078,15'd15398,15'd15718,15'd16038,15'd16358,15'd16678,15'd16998,15'd17318,15'd17638,15'd17958,15'd18278,15'd18598,15'd18918,15'd19238,15'd19558,15'd19878,15'd20198,15'd20518,15'd20838,15'd21158,15'd21478,15'd21798,15'd22118,15'd22438,15'd22758,15'd23078,15'd23398,15'd23718,15'd24038,15'd24358,15'd24678,15'd24998,15'd25318,
15'd37,15'd357,15'd677,15'd997,15'd1317,15'd1637,15'd1957,15'd2277,15'd2597,15'd2917,15'd3237,15'd3557,15'd3877,15'd4197,15'd4517,15'd4837,15'd5157,15'd5477,15'd5797,15'd6117,15'd6437,15'd6757,15'd7077,15'd7397,15'd7717,15'd8037,15'd8357,15'd8677,15'd8997,15'd9317,15'd9637,15'd9957,15'd10277,15'd10597,15'd10917,15'd11237,15'd11557,15'd11877,15'd12197,15'd12517,15'd12837,15'd13157,15'd13477,15'd13797,15'd14117,15'd14437,15'd14757,15'd15077,15'd15397,15'd15717,15'd16037,15'd16357,15'd16677,15'd16997,15'd17317,15'd17637,15'd17957,15'd18277,15'd18597,15'd18917,15'd19237,15'd19557,15'd19877,15'd20197,15'd20517,15'd20837,15'd21157,15'd21477,15'd21797,15'd22117,15'd22437,15'd22757,15'd23077,15'd23397,15'd23717,15'd24037,15'd24357,15'd24677,15'd24997,15'd25317,
15'd36,15'd356,15'd676,15'd996,15'd1316,15'd1636,15'd1956,15'd2276,15'd2596,15'd2916,15'd3236,15'd3556,15'd3876,15'd4196,15'd4516,15'd4836,15'd5156,15'd5476,15'd5796,15'd6116,15'd6436,15'd6756,15'd7076,15'd7396,15'd7716,15'd8036,15'd8356,15'd8676,15'd8996,15'd9316,15'd9636,15'd9956,15'd10276,15'd10596,15'd10916,15'd11236,15'd11556,15'd11876,15'd12196,15'd12516,15'd12836,15'd13156,15'd13476,15'd13796,15'd14116,15'd14436,15'd14756,15'd15076,15'd15396,15'd15716,15'd16036,15'd16356,15'd16676,15'd16996,15'd17316,15'd17636,15'd17956,15'd18276,15'd18596,15'd18916,15'd19236,15'd19556,15'd19876,15'd20196,15'd20516,15'd20836,15'd21156,15'd21476,15'd21796,15'd22116,15'd22436,15'd22756,15'd23076,15'd23396,15'd23716,15'd24036,15'd24356,15'd24676,15'd24996,15'd25316,
15'd35,15'd355,15'd675,15'd995,15'd1315,15'd1635,15'd1955,15'd2275,15'd2595,15'd2915,15'd3235,15'd3555,15'd3875,15'd4195,15'd4515,15'd4835,15'd5155,15'd5475,15'd5795,15'd6115,15'd6435,15'd6755,15'd7075,15'd7395,15'd7715,15'd8035,15'd8355,15'd8675,15'd8995,15'd9315,15'd9635,15'd9955,15'd10275,15'd10595,15'd10915,15'd11235,15'd11555,15'd11875,15'd12195,15'd12515,15'd12835,15'd13155,15'd13475,15'd13795,15'd14115,15'd14435,15'd14755,15'd15075,15'd15395,15'd15715,15'd16035,15'd16355,15'd16675,15'd16995,15'd17315,15'd17635,15'd17955,15'd18275,15'd18595,15'd18915,15'd19235,15'd19555,15'd19875,15'd20195,15'd20515,15'd20835,15'd21155,15'd21475,15'd21795,15'd22115,15'd22435,15'd22755,15'd23075,15'd23395,15'd23715,15'd24035,15'd24355,15'd24675,15'd24995,15'd25315,
15'd34,15'd354,15'd674,15'd994,15'd1314,15'd1634,15'd1954,15'd2274,15'd2594,15'd2914,15'd3234,15'd3554,15'd3874,15'd4194,15'd4514,15'd4834,15'd5154,15'd5474,15'd5794,15'd6114,15'd6434,15'd6754,15'd7074,15'd7394,15'd7714,15'd8034,15'd8354,15'd8674,15'd8994,15'd9314,15'd9634,15'd9954,15'd10274,15'd10594,15'd10914,15'd11234,15'd11554,15'd11874,15'd12194,15'd12514,15'd12834,15'd13154,15'd13474,15'd13794,15'd14114,15'd14434,15'd14754,15'd15074,15'd15394,15'd15714,15'd16034,15'd16354,15'd16674,15'd16994,15'd17314,15'd17634,15'd17954,15'd18274,15'd18594,15'd18914,15'd19234,15'd19554,15'd19874,15'd20194,15'd20514,15'd20834,15'd21154,15'd21474,15'd21794,15'd22114,15'd22434,15'd22754,15'd23074,15'd23394,15'd23714,15'd24034,15'd24354,15'd24674,15'd24994,15'd25314,
15'd33,15'd353,15'd673,15'd993,15'd1313,15'd1633,15'd1953,15'd2273,15'd2593,15'd2913,15'd3233,15'd3553,15'd3873,15'd4193,15'd4513,15'd4833,15'd5153,15'd5473,15'd5793,15'd6113,15'd6433,15'd6753,15'd7073,15'd7393,15'd7713,15'd8033,15'd8353,15'd8673,15'd8993,15'd9313,15'd9633,15'd9953,15'd10273,15'd10593,15'd10913,15'd11233,15'd11553,15'd11873,15'd12193,15'd12513,15'd12833,15'd13153,15'd13473,15'd13793,15'd14113,15'd14433,15'd14753,15'd15073,15'd15393,15'd15713,15'd16033,15'd16353,15'd16673,15'd16993,15'd17313,15'd17633,15'd17953,15'd18273,15'd18593,15'd18913,15'd19233,15'd19553,15'd19873,15'd20193,15'd20513,15'd20833,15'd21153,15'd21473,15'd21793,15'd22113,15'd22433,15'd22753,15'd23073,15'd23393,15'd23713,15'd24033,15'd24353,15'd24673,15'd24993,15'd25313,
15'd32,15'd352,15'd672,15'd992,15'd1312,15'd1632,15'd1952,15'd2272,15'd2592,15'd2912,15'd3232,15'd3552,15'd3872,15'd4192,15'd4512,15'd4832,15'd5152,15'd5472,15'd5792,15'd6112,15'd6432,15'd6752,15'd7072,15'd7392,15'd7712,15'd8032,15'd8352,15'd8672,15'd8992,15'd9312,15'd9632,15'd9952,15'd10272,15'd10592,15'd10912,15'd11232,15'd11552,15'd11872,15'd12192,15'd12512,15'd12832,15'd13152,15'd13472,15'd13792,15'd14112,15'd14432,15'd14752,15'd15072,15'd15392,15'd15712,15'd16032,15'd16352,15'd16672,15'd16992,15'd17312,15'd17632,15'd17952,15'd18272,15'd18592,15'd18912,15'd19232,15'd19552,15'd19872,15'd20192,15'd20512,15'd20832,15'd21152,15'd21472,15'd21792,15'd22112,15'd22432,15'd22752,15'd23072,15'd23392,15'd23712,15'd24032,15'd24352,15'd24672,15'd24992,15'd25312,
15'd31,15'd351,15'd671,15'd991,15'd1311,15'd1631,15'd1951,15'd2271,15'd2591,15'd2911,15'd3231,15'd3551,15'd3871,15'd4191,15'd4511,15'd4831,15'd5151,15'd5471,15'd5791,15'd6111,15'd6431,15'd6751,15'd7071,15'd7391,15'd7711,15'd8031,15'd8351,15'd8671,15'd8991,15'd9311,15'd9631,15'd9951,15'd10271,15'd10591,15'd10911,15'd11231,15'd11551,15'd11871,15'd12191,15'd12511,15'd12831,15'd13151,15'd13471,15'd13791,15'd14111,15'd14431,15'd14751,15'd15071,15'd15391,15'd15711,15'd16031,15'd16351,15'd16671,15'd16991,15'd17311,15'd17631,15'd17951,15'd18271,15'd18591,15'd18911,15'd19231,15'd19551,15'd19871,15'd20191,15'd20511,15'd20831,15'd21151,15'd21471,15'd21791,15'd22111,15'd22431,15'd22751,15'd23071,15'd23391,15'd23711,15'd24031,15'd24351,15'd24671,15'd24991,15'd25311,
15'd30,15'd350,15'd670,15'd990,15'd1310,15'd1630,15'd1950,15'd2270,15'd2590,15'd2910,15'd3230,15'd3550,15'd3870,15'd4190,15'd4510,15'd4830,15'd5150,15'd5470,15'd5790,15'd6110,15'd6430,15'd6750,15'd7070,15'd7390,15'd7710,15'd8030,15'd8350,15'd8670,15'd8990,15'd9310,15'd9630,15'd9950,15'd10270,15'd10590,15'd10910,15'd11230,15'd11550,15'd11870,15'd12190,15'd12510,15'd12830,15'd13150,15'd13470,15'd13790,15'd14110,15'd14430,15'd14750,15'd15070,15'd15390,15'd15710,15'd16030,15'd16350,15'd16670,15'd16990,15'd17310,15'd17630,15'd17950,15'd18270,15'd18590,15'd18910,15'd19230,15'd19550,15'd19870,15'd20190,15'd20510,15'd20830,15'd21150,15'd21470,15'd21790,15'd22110,15'd22430,15'd22750,15'd23070,15'd23390,15'd23710,15'd24030,15'd24350,15'd24670,15'd24990,15'd25310,
15'd29,15'd349,15'd669,15'd989,15'd1309,15'd1629,15'd1949,15'd2269,15'd2589,15'd2909,15'd3229,15'd3549,15'd3869,15'd4189,15'd4509,15'd4829,15'd5149,15'd5469,15'd5789,15'd6109,15'd6429,15'd6749,15'd7069,15'd7389,15'd7709,15'd8029,15'd8349,15'd8669,15'd8989,15'd9309,15'd9629,15'd9949,15'd10269,15'd10589,15'd10909,15'd11229,15'd11549,15'd11869,15'd12189,15'd12509,15'd12829,15'd13149,15'd13469,15'd13789,15'd14109,15'd14429,15'd14749,15'd15069,15'd15389,15'd15709,15'd16029,15'd16349,15'd16669,15'd16989,15'd17309,15'd17629,15'd17949,15'd18269,15'd18589,15'd18909,15'd19229,15'd19549,15'd19869,15'd20189,15'd20509,15'd20829,15'd21149,15'd21469,15'd21789,15'd22109,15'd22429,15'd22749,15'd23069,15'd23389,15'd23709,15'd24029,15'd24349,15'd24669,15'd24989,15'd25309,
15'd28,15'd348,15'd668,15'd988,15'd1308,15'd1628,15'd1948,15'd2268,15'd2588,15'd2908,15'd3228,15'd3548,15'd3868,15'd4188,15'd4508,15'd4828,15'd5148,15'd5468,15'd5788,15'd6108,15'd6428,15'd6748,15'd7068,15'd7388,15'd7708,15'd8028,15'd8348,15'd8668,15'd8988,15'd9308,15'd9628,15'd9948,15'd10268,15'd10588,15'd10908,15'd11228,15'd11548,15'd11868,15'd12188,15'd12508,15'd12828,15'd13148,15'd13468,15'd13788,15'd14108,15'd14428,15'd14748,15'd15068,15'd15388,15'd15708,15'd16028,15'd16348,15'd16668,15'd16988,15'd17308,15'd17628,15'd17948,15'd18268,15'd18588,15'd18908,15'd19228,15'd19548,15'd19868,15'd20188,15'd20508,15'd20828,15'd21148,15'd21468,15'd21788,15'd22108,15'd22428,15'd22748,15'd23068,15'd23388,15'd23708,15'd24028,15'd24348,15'd24668,15'd24988,15'd25308,
15'd27,15'd347,15'd667,15'd987,15'd1307,15'd1627,15'd1947,15'd2267,15'd2587,15'd2907,15'd3227,15'd3547,15'd3867,15'd4187,15'd4507,15'd4827,15'd5147,15'd5467,15'd5787,15'd6107,15'd6427,15'd6747,15'd7067,15'd7387,15'd7707,15'd8027,15'd8347,15'd8667,15'd8987,15'd9307,15'd9627,15'd9947,15'd10267,15'd10587,15'd10907,15'd11227,15'd11547,15'd11867,15'd12187,15'd12507,15'd12827,15'd13147,15'd13467,15'd13787,15'd14107,15'd14427,15'd14747,15'd15067,15'd15387,15'd15707,15'd16027,15'd16347,15'd16667,15'd16987,15'd17307,15'd17627,15'd17947,15'd18267,15'd18587,15'd18907,15'd19227,15'd19547,15'd19867,15'd20187,15'd20507,15'd20827,15'd21147,15'd21467,15'd21787,15'd22107,15'd22427,15'd22747,15'd23067,15'd23387,15'd23707,15'd24027,15'd24347,15'd24667,15'd24987,15'd25307,
15'd26,15'd346,15'd666,15'd986,15'd1306,15'd1626,15'd1946,15'd2266,15'd2586,15'd2906,15'd3226,15'd3546,15'd3866,15'd4186,15'd4506,15'd4826,15'd5146,15'd5466,15'd5786,15'd6106,15'd6426,15'd6746,15'd7066,15'd7386,15'd7706,15'd8026,15'd8346,15'd8666,15'd8986,15'd9306,15'd9626,15'd9946,15'd10266,15'd10586,15'd10906,15'd11226,15'd11546,15'd11866,15'd12186,15'd12506,15'd12826,15'd13146,15'd13466,15'd13786,15'd14106,15'd14426,15'd14746,15'd15066,15'd15386,15'd15706,15'd16026,15'd16346,15'd16666,15'd16986,15'd17306,15'd17626,15'd17946,15'd18266,15'd18586,15'd18906,15'd19226,15'd19546,15'd19866,15'd20186,15'd20506,15'd20826,15'd21146,15'd21466,15'd21786,15'd22106,15'd22426,15'd22746,15'd23066,15'd23386,15'd23706,15'd24026,15'd24346,15'd24666,15'd24986,15'd25306,
15'd25,15'd345,15'd665,15'd985,15'd1305,15'd1625,15'd1945,15'd2265,15'd2585,15'd2905,15'd3225,15'd3545,15'd3865,15'd4185,15'd4505,15'd4825,15'd5145,15'd5465,15'd5785,15'd6105,15'd6425,15'd6745,15'd7065,15'd7385,15'd7705,15'd8025,15'd8345,15'd8665,15'd8985,15'd9305,15'd9625,15'd9945,15'd10265,15'd10585,15'd10905,15'd11225,15'd11545,15'd11865,15'd12185,15'd12505,15'd12825,15'd13145,15'd13465,15'd13785,15'd14105,15'd14425,15'd14745,15'd15065,15'd15385,15'd15705,15'd16025,15'd16345,15'd16665,15'd16985,15'd17305,15'd17625,15'd17945,15'd18265,15'd18585,15'd18905,15'd19225,15'd19545,15'd19865,15'd20185,15'd20505,15'd20825,15'd21145,15'd21465,15'd21785,15'd22105,15'd22425,15'd22745,15'd23065,15'd23385,15'd23705,15'd24025,15'd24345,15'd24665,15'd24985,15'd25305,
15'd24,15'd344,15'd664,15'd984,15'd1304,15'd1624,15'd1944,15'd2264,15'd2584,15'd2904,15'd3224,15'd3544,15'd3864,15'd4184,15'd4504,15'd4824,15'd5144,15'd5464,15'd5784,15'd6104,15'd6424,15'd6744,15'd7064,15'd7384,15'd7704,15'd8024,15'd8344,15'd8664,15'd8984,15'd9304,15'd9624,15'd9944,15'd10264,15'd10584,15'd10904,15'd11224,15'd11544,15'd11864,15'd12184,15'd12504,15'd12824,15'd13144,15'd13464,15'd13784,15'd14104,15'd14424,15'd14744,15'd15064,15'd15384,15'd15704,15'd16024,15'd16344,15'd16664,15'd16984,15'd17304,15'd17624,15'd17944,15'd18264,15'd18584,15'd18904,15'd19224,15'd19544,15'd19864,15'd20184,15'd20504,15'd20824,15'd21144,15'd21464,15'd21784,15'd22104,15'd22424,15'd22744,15'd23064,15'd23384,15'd23704,15'd24024,15'd24344,15'd24664,15'd24984,15'd25304,
15'd23,15'd343,15'd663,15'd983,15'd1303,15'd1623,15'd1943,15'd2263,15'd2583,15'd2903,15'd3223,15'd3543,15'd3863,15'd4183,15'd4503,15'd4823,15'd5143,15'd5463,15'd5783,15'd6103,15'd6423,15'd6743,15'd7063,15'd7383,15'd7703,15'd8023,15'd8343,15'd8663,15'd8983,15'd9303,15'd9623,15'd9943,15'd10263,15'd10583,15'd10903,15'd11223,15'd11543,15'd11863,15'd12183,15'd12503,15'd12823,15'd13143,15'd13463,15'd13783,15'd14103,15'd14423,15'd14743,15'd15063,15'd15383,15'd15703,15'd16023,15'd16343,15'd16663,15'd16983,15'd17303,15'd17623,15'd17943,15'd18263,15'd18583,15'd18903,15'd19223,15'd19543,15'd19863,15'd20183,15'd20503,15'd20823,15'd21143,15'd21463,15'd21783,15'd22103,15'd22423,15'd22743,15'd23063,15'd23383,15'd23703,15'd24023,15'd24343,15'd24663,15'd24983,15'd25303,
15'd22,15'd342,15'd662,15'd982,15'd1302,15'd1622,15'd1942,15'd2262,15'd2582,15'd2902,15'd3222,15'd3542,15'd3862,15'd4182,15'd4502,15'd4822,15'd5142,15'd5462,15'd5782,15'd6102,15'd6422,15'd6742,15'd7062,15'd7382,15'd7702,15'd8022,15'd8342,15'd8662,15'd8982,15'd9302,15'd9622,15'd9942,15'd10262,15'd10582,15'd10902,15'd11222,15'd11542,15'd11862,15'd12182,15'd12502,15'd12822,15'd13142,15'd13462,15'd13782,15'd14102,15'd14422,15'd14742,15'd15062,15'd15382,15'd15702,15'd16022,15'd16342,15'd16662,15'd16982,15'd17302,15'd17622,15'd17942,15'd18262,15'd18582,15'd18902,15'd19222,15'd19542,15'd19862,15'd20182,15'd20502,15'd20822,15'd21142,15'd21462,15'd21782,15'd22102,15'd22422,15'd22742,15'd23062,15'd23382,15'd23702,15'd24022,15'd24342,15'd24662,15'd24982,15'd25302,
15'd21,15'd341,15'd661,15'd981,15'd1301,15'd1621,15'd1941,15'd2261,15'd2581,15'd2901,15'd3221,15'd3541,15'd3861,15'd4181,15'd4501,15'd4821,15'd5141,15'd5461,15'd5781,15'd6101,15'd6421,15'd6741,15'd7061,15'd7381,15'd7701,15'd8021,15'd8341,15'd8661,15'd8981,15'd9301,15'd9621,15'd9941,15'd10261,15'd10581,15'd10901,15'd11221,15'd11541,15'd11861,15'd12181,15'd12501,15'd12821,15'd13141,15'd13461,15'd13781,15'd14101,15'd14421,15'd14741,15'd15061,15'd15381,15'd15701,15'd16021,15'd16341,15'd16661,15'd16981,15'd17301,15'd17621,15'd17941,15'd18261,15'd18581,15'd18901,15'd19221,15'd19541,15'd19861,15'd20181,15'd20501,15'd20821,15'd21141,15'd21461,15'd21781,15'd22101,15'd22421,15'd22741,15'd23061,15'd23381,15'd23701,15'd24021,15'd24341,15'd24661,15'd24981,15'd25301,
15'd20,15'd340,15'd660,15'd980,15'd1300,15'd1620,15'd1940,15'd2260,15'd2580,15'd2900,15'd3220,15'd3540,15'd3860,15'd4180,15'd4500,15'd4820,15'd5140,15'd5460,15'd5780,15'd6100,15'd6420,15'd6740,15'd7060,15'd7380,15'd7700,15'd8020,15'd8340,15'd8660,15'd8980,15'd9300,15'd9620,15'd9940,15'd10260,15'd10580,15'd10900,15'd11220,15'd11540,15'd11860,15'd12180,15'd12500,15'd12820,15'd13140,15'd13460,15'd13780,15'd14100,15'd14420,15'd14740,15'd15060,15'd15380,15'd15700,15'd16020,15'd16340,15'd16660,15'd16980,15'd17300,15'd17620,15'd17940,15'd18260,15'd18580,15'd18900,15'd19220,15'd19540,15'd19860,15'd20180,15'd20500,15'd20820,15'd21140,15'd21460,15'd21780,15'd22100,15'd22420,15'd22740,15'd23060,15'd23380,15'd23700,15'd24020,15'd24340,15'd24660,15'd24980,15'd25300,
15'd19,15'd339,15'd659,15'd979,15'd1299,15'd1619,15'd1939,15'd2259,15'd2579,15'd2899,15'd3219,15'd3539,15'd3859,15'd4179,15'd4499,15'd4819,15'd5139,15'd5459,15'd5779,15'd6099,15'd6419,15'd6739,15'd7059,15'd7379,15'd7699,15'd8019,15'd8339,15'd8659,15'd8979,15'd9299,15'd9619,15'd9939,15'd10259,15'd10579,15'd10899,15'd11219,15'd11539,15'd11859,15'd12179,15'd12499,15'd12819,15'd13139,15'd13459,15'd13779,15'd14099,15'd14419,15'd14739,15'd15059,15'd15379,15'd15699,15'd16019,15'd16339,15'd16659,15'd16979,15'd17299,15'd17619,15'd17939,15'd18259,15'd18579,15'd18899,15'd19219,15'd19539,15'd19859,15'd20179,15'd20499,15'd20819,15'd21139,15'd21459,15'd21779,15'd22099,15'd22419,15'd22739,15'd23059,15'd23379,15'd23699,15'd24019,15'd24339,15'd24659,15'd24979,15'd25299,
15'd18,15'd338,15'd658,15'd978,15'd1298,15'd1618,15'd1938,15'd2258,15'd2578,15'd2898,15'd3218,15'd3538,15'd3858,15'd4178,15'd4498,15'd4818,15'd5138,15'd5458,15'd5778,15'd6098,15'd6418,15'd6738,15'd7058,15'd7378,15'd7698,15'd8018,15'd8338,15'd8658,15'd8978,15'd9298,15'd9618,15'd9938,15'd10258,15'd10578,15'd10898,15'd11218,15'd11538,15'd11858,15'd12178,15'd12498,15'd12818,15'd13138,15'd13458,15'd13778,15'd14098,15'd14418,15'd14738,15'd15058,15'd15378,15'd15698,15'd16018,15'd16338,15'd16658,15'd16978,15'd17298,15'd17618,15'd17938,15'd18258,15'd18578,15'd18898,15'd19218,15'd19538,15'd19858,15'd20178,15'd20498,15'd20818,15'd21138,15'd21458,15'd21778,15'd22098,15'd22418,15'd22738,15'd23058,15'd23378,15'd23698,15'd24018,15'd24338,15'd24658,15'd24978,15'd25298,
15'd17,15'd337,15'd657,15'd977,15'd1297,15'd1617,15'd1937,15'd2257,15'd2577,15'd2897,15'd3217,15'd3537,15'd3857,15'd4177,15'd4497,15'd4817,15'd5137,15'd5457,15'd5777,15'd6097,15'd6417,15'd6737,15'd7057,15'd7377,15'd7697,15'd8017,15'd8337,15'd8657,15'd8977,15'd9297,15'd9617,15'd9937,15'd10257,15'd10577,15'd10897,15'd11217,15'd11537,15'd11857,15'd12177,15'd12497,15'd12817,15'd13137,15'd13457,15'd13777,15'd14097,15'd14417,15'd14737,15'd15057,15'd15377,15'd15697,15'd16017,15'd16337,15'd16657,15'd16977,15'd17297,15'd17617,15'd17937,15'd18257,15'd18577,15'd18897,15'd19217,15'd19537,15'd19857,15'd20177,15'd20497,15'd20817,15'd21137,15'd21457,15'd21777,15'd22097,15'd22417,15'd22737,15'd23057,15'd23377,15'd23697,15'd24017,15'd24337,15'd24657,15'd24977,15'd25297,
15'd16,15'd336,15'd656,15'd976,15'd1296,15'd1616,15'd1936,15'd2256,15'd2576,15'd2896,15'd3216,15'd3536,15'd3856,15'd4176,15'd4496,15'd4816,15'd5136,15'd5456,15'd5776,15'd6096,15'd6416,15'd6736,15'd7056,15'd7376,15'd7696,15'd8016,15'd8336,15'd8656,15'd8976,15'd9296,15'd9616,15'd9936,15'd10256,15'd10576,15'd10896,15'd11216,15'd11536,15'd11856,15'd12176,15'd12496,15'd12816,15'd13136,15'd13456,15'd13776,15'd14096,15'd14416,15'd14736,15'd15056,15'd15376,15'd15696,15'd16016,15'd16336,15'd16656,15'd16976,15'd17296,15'd17616,15'd17936,15'd18256,15'd18576,15'd18896,15'd19216,15'd19536,15'd19856,15'd20176,15'd20496,15'd20816,15'd21136,15'd21456,15'd21776,15'd22096,15'd22416,15'd22736,15'd23056,15'd23376,15'd23696,15'd24016,15'd24336,15'd24656,15'd24976,15'd25296,
15'd15,15'd335,15'd655,15'd975,15'd1295,15'd1615,15'd1935,15'd2255,15'd2575,15'd2895,15'd3215,15'd3535,15'd3855,15'd4175,15'd4495,15'd4815,15'd5135,15'd5455,15'd5775,15'd6095,15'd6415,15'd6735,15'd7055,15'd7375,15'd7695,15'd8015,15'd8335,15'd8655,15'd8975,15'd9295,15'd9615,15'd9935,15'd10255,15'd10575,15'd10895,15'd11215,15'd11535,15'd11855,15'd12175,15'd12495,15'd12815,15'd13135,15'd13455,15'd13775,15'd14095,15'd14415,15'd14735,15'd15055,15'd15375,15'd15695,15'd16015,15'd16335,15'd16655,15'd16975,15'd17295,15'd17615,15'd17935,15'd18255,15'd18575,15'd18895,15'd19215,15'd19535,15'd19855,15'd20175,15'd20495,15'd20815,15'd21135,15'd21455,15'd21775,15'd22095,15'd22415,15'd22735,15'd23055,15'd23375,15'd23695,15'd24015,15'd24335,15'd24655,15'd24975,15'd25295,
15'd14,15'd334,15'd654,15'd974,15'd1294,15'd1614,15'd1934,15'd2254,15'd2574,15'd2894,15'd3214,15'd3534,15'd3854,15'd4174,15'd4494,15'd4814,15'd5134,15'd5454,15'd5774,15'd6094,15'd6414,15'd6734,15'd7054,15'd7374,15'd7694,15'd8014,15'd8334,15'd8654,15'd8974,15'd9294,15'd9614,15'd9934,15'd10254,15'd10574,15'd10894,15'd11214,15'd11534,15'd11854,15'd12174,15'd12494,15'd12814,15'd13134,15'd13454,15'd13774,15'd14094,15'd14414,15'd14734,15'd15054,15'd15374,15'd15694,15'd16014,15'd16334,15'd16654,15'd16974,15'd17294,15'd17614,15'd17934,15'd18254,15'd18574,15'd18894,15'd19214,15'd19534,15'd19854,15'd20174,15'd20494,15'd20814,15'd21134,15'd21454,15'd21774,15'd22094,15'd22414,15'd22734,15'd23054,15'd23374,15'd23694,15'd24014,15'd24334,15'd24654,15'd24974,15'd25294,
15'd13,15'd333,15'd653,15'd973,15'd1293,15'd1613,15'd1933,15'd2253,15'd2573,15'd2893,15'd3213,15'd3533,15'd3853,15'd4173,15'd4493,15'd4813,15'd5133,15'd5453,15'd5773,15'd6093,15'd6413,15'd6733,15'd7053,15'd7373,15'd7693,15'd8013,15'd8333,15'd8653,15'd8973,15'd9293,15'd9613,15'd9933,15'd10253,15'd10573,15'd10893,15'd11213,15'd11533,15'd11853,15'd12173,15'd12493,15'd12813,15'd13133,15'd13453,15'd13773,15'd14093,15'd14413,15'd14733,15'd15053,15'd15373,15'd15693,15'd16013,15'd16333,15'd16653,15'd16973,15'd17293,15'd17613,15'd17933,15'd18253,15'd18573,15'd18893,15'd19213,15'd19533,15'd19853,15'd20173,15'd20493,15'd20813,15'd21133,15'd21453,15'd21773,15'd22093,15'd22413,15'd22733,15'd23053,15'd23373,15'd23693,15'd24013,15'd24333,15'd24653,15'd24973,15'd25293,
15'd12,15'd332,15'd652,15'd972,15'd1292,15'd1612,15'd1932,15'd2252,15'd2572,15'd2892,15'd3212,15'd3532,15'd3852,15'd4172,15'd4492,15'd4812,15'd5132,15'd5452,15'd5772,15'd6092,15'd6412,15'd6732,15'd7052,15'd7372,15'd7692,15'd8012,15'd8332,15'd8652,15'd8972,15'd9292,15'd9612,15'd9932,15'd10252,15'd10572,15'd10892,15'd11212,15'd11532,15'd11852,15'd12172,15'd12492,15'd12812,15'd13132,15'd13452,15'd13772,15'd14092,15'd14412,15'd14732,15'd15052,15'd15372,15'd15692,15'd16012,15'd16332,15'd16652,15'd16972,15'd17292,15'd17612,15'd17932,15'd18252,15'd18572,15'd18892,15'd19212,15'd19532,15'd19852,15'd20172,15'd20492,15'd20812,15'd21132,15'd21452,15'd21772,15'd22092,15'd22412,15'd22732,15'd23052,15'd23372,15'd23692,15'd24012,15'd24332,15'd24652,15'd24972,15'd25292,
15'd11,15'd331,15'd651,15'd971,15'd1291,15'd1611,15'd1931,15'd2251,15'd2571,15'd2891,15'd3211,15'd3531,15'd3851,15'd4171,15'd4491,15'd4811,15'd5131,15'd5451,15'd5771,15'd6091,15'd6411,15'd6731,15'd7051,15'd7371,15'd7691,15'd8011,15'd8331,15'd8651,15'd8971,15'd9291,15'd9611,15'd9931,15'd10251,15'd10571,15'd10891,15'd11211,15'd11531,15'd11851,15'd12171,15'd12491,15'd12811,15'd13131,15'd13451,15'd13771,15'd14091,15'd14411,15'd14731,15'd15051,15'd15371,15'd15691,15'd16011,15'd16331,15'd16651,15'd16971,15'd17291,15'd17611,15'd17931,15'd18251,15'd18571,15'd18891,15'd19211,15'd19531,15'd19851,15'd20171,15'd20491,15'd20811,15'd21131,15'd21451,15'd21771,15'd22091,15'd22411,15'd22731,15'd23051,15'd23371,15'd23691,15'd24011,15'd24331,15'd24651,15'd24971,15'd25291,
15'd10,15'd330,15'd650,15'd970,15'd1290,15'd1610,15'd1930,15'd2250,15'd2570,15'd2890,15'd3210,15'd3530,15'd3850,15'd4170,15'd4490,15'd4810,15'd5130,15'd5450,15'd5770,15'd6090,15'd6410,15'd6730,15'd7050,15'd7370,15'd7690,15'd8010,15'd8330,15'd8650,15'd8970,15'd9290,15'd9610,15'd9930,15'd10250,15'd10570,15'd10890,15'd11210,15'd11530,15'd11850,15'd12170,15'd12490,15'd12810,15'd13130,15'd13450,15'd13770,15'd14090,15'd14410,15'd14730,15'd15050,15'd15370,15'd15690,15'd16010,15'd16330,15'd16650,15'd16970,15'd17290,15'd17610,15'd17930,15'd18250,15'd18570,15'd18890,15'd19210,15'd19530,15'd19850,15'd20170,15'd20490,15'd20810,15'd21130,15'd21450,15'd21770,15'd22090,15'd22410,15'd22730,15'd23050,15'd23370,15'd23690,15'd24010,15'd24330,15'd24650,15'd24970,15'd25290,
15'd9,15'd329,15'd649,15'd969,15'd1289,15'd1609,15'd1929,15'd2249,15'd2569,15'd2889,15'd3209,15'd3529,15'd3849,15'd4169,15'd4489,15'd4809,15'd5129,15'd5449,15'd5769,15'd6089,15'd6409,15'd6729,15'd7049,15'd7369,15'd7689,15'd8009,15'd8329,15'd8649,15'd8969,15'd9289,15'd9609,15'd9929,15'd10249,15'd10569,15'd10889,15'd11209,15'd11529,15'd11849,15'd12169,15'd12489,15'd12809,15'd13129,15'd13449,15'd13769,15'd14089,15'd14409,15'd14729,15'd15049,15'd15369,15'd15689,15'd16009,15'd16329,15'd16649,15'd16969,15'd17289,15'd17609,15'd17929,15'd18249,15'd18569,15'd18889,15'd19209,15'd19529,15'd19849,15'd20169,15'd20489,15'd20809,15'd21129,15'd21449,15'd21769,15'd22089,15'd22409,15'd22729,15'd23049,15'd23369,15'd23689,15'd24009,15'd24329,15'd24649,15'd24969,15'd25289,
15'd8,15'd328,15'd648,15'd968,15'd1288,15'd1608,15'd1928,15'd2248,15'd2568,15'd2888,15'd3208,15'd3528,15'd3848,15'd4168,15'd4488,15'd4808,15'd5128,15'd5448,15'd5768,15'd6088,15'd6408,15'd6728,15'd7048,15'd7368,15'd7688,15'd8008,15'd8328,15'd8648,15'd8968,15'd9288,15'd9608,15'd9928,15'd10248,15'd10568,15'd10888,15'd11208,15'd11528,15'd11848,15'd12168,15'd12488,15'd12808,15'd13128,15'd13448,15'd13768,15'd14088,15'd14408,15'd14728,15'd15048,15'd15368,15'd15688,15'd16008,15'd16328,15'd16648,15'd16968,15'd17288,15'd17608,15'd17928,15'd18248,15'd18568,15'd18888,15'd19208,15'd19528,15'd19848,15'd20168,15'd20488,15'd20808,15'd21128,15'd21448,15'd21768,15'd22088,15'd22408,15'd22728,15'd23048,15'd23368,15'd23688,15'd24008,15'd24328,15'd24648,15'd24968,15'd25288,
15'd7,15'd327,15'd647,15'd967,15'd1287,15'd1607,15'd1927,15'd2247,15'd2567,15'd2887,15'd3207,15'd3527,15'd3847,15'd4167,15'd4487,15'd4807,15'd5127,15'd5447,15'd5767,15'd6087,15'd6407,15'd6727,15'd7047,15'd7367,15'd7687,15'd8007,15'd8327,15'd8647,15'd8967,15'd9287,15'd9607,15'd9927,15'd10247,15'd10567,15'd10887,15'd11207,15'd11527,15'd11847,15'd12167,15'd12487,15'd12807,15'd13127,15'd13447,15'd13767,15'd14087,15'd14407,15'd14727,15'd15047,15'd15367,15'd15687,15'd16007,15'd16327,15'd16647,15'd16967,15'd17287,15'd17607,15'd17927,15'd18247,15'd18567,15'd18887,15'd19207,15'd19527,15'd19847,15'd20167,15'd20487,15'd20807,15'd21127,15'd21447,15'd21767,15'd22087,15'd22407,15'd22727,15'd23047,15'd23367,15'd23687,15'd24007,15'd24327,15'd24647,15'd24967,15'd25287,
15'd6,15'd326,15'd646,15'd966,15'd1286,15'd1606,15'd1926,15'd2246,15'd2566,15'd2886,15'd3206,15'd3526,15'd3846,15'd4166,15'd4486,15'd4806,15'd5126,15'd5446,15'd5766,15'd6086,15'd6406,15'd6726,15'd7046,15'd7366,15'd7686,15'd8006,15'd8326,15'd8646,15'd8966,15'd9286,15'd9606,15'd9926,15'd10246,15'd10566,15'd10886,15'd11206,15'd11526,15'd11846,15'd12166,15'd12486,15'd12806,15'd13126,15'd13446,15'd13766,15'd14086,15'd14406,15'd14726,15'd15046,15'd15366,15'd15686,15'd16006,15'd16326,15'd16646,15'd16966,15'd17286,15'd17606,15'd17926,15'd18246,15'd18566,15'd18886,15'd19206,15'd19526,15'd19846,15'd20166,15'd20486,15'd20806,15'd21126,15'd21446,15'd21766,15'd22086,15'd22406,15'd22726,15'd23046,15'd23366,15'd23686,15'd24006,15'd24326,15'd24646,15'd24966,15'd25286,
15'd5,15'd325,15'd645,15'd965,15'd1285,15'd1605,15'd1925,15'd2245,15'd2565,15'd2885,15'd3205,15'd3525,15'd3845,15'd4165,15'd4485,15'd4805,15'd5125,15'd5445,15'd5765,15'd6085,15'd6405,15'd6725,15'd7045,15'd7365,15'd7685,15'd8005,15'd8325,15'd8645,15'd8965,15'd9285,15'd9605,15'd9925,15'd10245,15'd10565,15'd10885,15'd11205,15'd11525,15'd11845,15'd12165,15'd12485,15'd12805,15'd13125,15'd13445,15'd13765,15'd14085,15'd14405,15'd14725,15'd15045,15'd15365,15'd15685,15'd16005,15'd16325,15'd16645,15'd16965,15'd17285,15'd17605,15'd17925,15'd18245,15'd18565,15'd18885,15'd19205,15'd19525,15'd19845,15'd20165,15'd20485,15'd20805,15'd21125,15'd21445,15'd21765,15'd22085,15'd22405,15'd22725,15'd23045,15'd23365,15'd23685,15'd24005,15'd24325,15'd24645,15'd24965,15'd25285,
15'd4,15'd324,15'd644,15'd964,15'd1284,15'd1604,15'd1924,15'd2244,15'd2564,15'd2884,15'd3204,15'd3524,15'd3844,15'd4164,15'd4484,15'd4804,15'd5124,15'd5444,15'd5764,15'd6084,15'd6404,15'd6724,15'd7044,15'd7364,15'd7684,15'd8004,15'd8324,15'd8644,15'd8964,15'd9284,15'd9604,15'd9924,15'd10244,15'd10564,15'd10884,15'd11204,15'd11524,15'd11844,15'd12164,15'd12484,15'd12804,15'd13124,15'd13444,15'd13764,15'd14084,15'd14404,15'd14724,15'd15044,15'd15364,15'd15684,15'd16004,15'd16324,15'd16644,15'd16964,15'd17284,15'd17604,15'd17924,15'd18244,15'd18564,15'd18884,15'd19204,15'd19524,15'd19844,15'd20164,15'd20484,15'd20804,15'd21124,15'd21444,15'd21764,15'd22084,15'd22404,15'd22724,15'd23044,15'd23364,15'd23684,15'd24004,15'd24324,15'd24644,15'd24964,15'd25284,
15'd3,15'd323,15'd643,15'd963,15'd1283,15'd1603,15'd1923,15'd2243,15'd2563,15'd2883,15'd3203,15'd3523,15'd3843,15'd4163,15'd4483,15'd4803,15'd5123,15'd5443,15'd5763,15'd6083,15'd6403,15'd6723,15'd7043,15'd7363,15'd7683,15'd8003,15'd8323,15'd8643,15'd8963,15'd9283,15'd9603,15'd9923,15'd10243,15'd10563,15'd10883,15'd11203,15'd11523,15'd11843,15'd12163,15'd12483,15'd12803,15'd13123,15'd13443,15'd13763,15'd14083,15'd14403,15'd14723,15'd15043,15'd15363,15'd15683,15'd16003,15'd16323,15'd16643,15'd16963,15'd17283,15'd17603,15'd17923,15'd18243,15'd18563,15'd18883,15'd19203,15'd19523,15'd19843,15'd20163,15'd20483,15'd20803,15'd21123,15'd21443,15'd21763,15'd22083,15'd22403,15'd22723,15'd23043,15'd23363,15'd23683,15'd24003,15'd24323,15'd24643,15'd24963,15'd25283,
15'd2,15'd322,15'd642,15'd962,15'd1282,15'd1602,15'd1922,15'd2242,15'd2562,15'd2882,15'd3202,15'd3522,15'd3842,15'd4162,15'd4482,15'd4802,15'd5122,15'd5442,15'd5762,15'd6082,15'd6402,15'd6722,15'd7042,15'd7362,15'd7682,15'd8002,15'd8322,15'd8642,15'd8962,15'd9282,15'd9602,15'd9922,15'd10242,15'd10562,15'd10882,15'd11202,15'd11522,15'd11842,15'd12162,15'd12482,15'd12802,15'd13122,15'd13442,15'd13762,15'd14082,15'd14402,15'd14722,15'd15042,15'd15362,15'd15682,15'd16002,15'd16322,15'd16642,15'd16962,15'd17282,15'd17602,15'd17922,15'd18242,15'd18562,15'd18882,15'd19202,15'd19522,15'd19842,15'd20162,15'd20482,15'd20802,15'd21122,15'd21442,15'd21762,15'd22082,15'd22402,15'd22722,15'd23042,15'd23362,15'd23682,15'd24002,15'd24322,15'd24642,15'd24962,15'd25282,
15'd1,15'd321,15'd641,15'd961,15'd1281,15'd1601,15'd1921,15'd2241,15'd2561,15'd2881,15'd3201,15'd3521,15'd3841,15'd4161,15'd4481,15'd4801,15'd5121,15'd5441,15'd5761,15'd6081,15'd6401,15'd6721,15'd7041,15'd7361,15'd7681,15'd8001,15'd8321,15'd8641,15'd8961,15'd9281,15'd9601,15'd9921,15'd10241,15'd10561,15'd10881,15'd11201,15'd11521,15'd11841,15'd12161,15'd12481,15'd12801,15'd13121,15'd13441,15'd13761,15'd14081,15'd14401,15'd14721,15'd15041,15'd15361,15'd15681,15'd16001,15'd16321,15'd16641,15'd16961,15'd17281,15'd17601,15'd17921,15'd18241,15'd18561,15'd18881,15'd19201,15'd19521,15'd19841,15'd20161,15'd20481,15'd20801,15'd21121,15'd21441,15'd21761,15'd22081,15'd22401,15'd22721,15'd23041,15'd23361,15'd23681,15'd24001,15'd24321,15'd24641,15'd24961,15'd25281,
15'd0,15'd320,15'd640,15'd960,15'd1280,15'd1600,15'd1920,15'd2240,15'd2560,15'd2880,15'd3200,15'd3520,15'd3840,15'd4160,15'd4480,15'd4800,15'd5120,15'd5440,15'd5760,15'd6080,15'd6400,15'd6720,15'd7040,15'd7360,15'd7680,15'd8000,15'd8320,15'd8640,15'd8960,15'd9280,15'd9600,15'd9920,15'd10240,15'd10560,15'd10880,15'd11200,15'd11520,15'd11840,15'd12160,15'd12480,15'd12800,15'd13120,15'd13440,15'd13760,15'd14080,15'd14400,15'd14720,15'd15040,15'd15360,15'd15680,15'd16000,15'd16320,15'd16640,15'd16960,15'd17280,15'd17600,15'd17920,15'd18240,15'd18560,15'd18880,15'd19200,15'd19520,15'd19840,15'd20160,15'd20480,15'd20800,15'd21120,15'd21440,15'd21760,15'd22080,15'd22400,15'd22720,15'd23040,15'd23360,15'd23680,15'd24000,15'd24320,15'd24640,15'd24960,15'd25280};
   
   
   
   assign pass = (zero==0 && one==0 && two==0 && three==0 && four==0 && five==0 && six==0 && seven==0 && eight==0 && nine==0 && ten==0 && ele==0) ? 1'b1 : 1'b0;

   always @ (posedge clk) begin
       
            if(hold == 1'b1) begin
                if( (h_cnt>>1)+320*(v_cnt>>1) < 25600 ) begin
                    if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 0 ) begin
                        pixel_addr <= state_0[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)) /320)*80 ];
                    end
                    else if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 1 ) begin
                        pixel_addr <= state_0[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)-80) /320)*80 ]+80;
                    end
                    else if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 2 ) begin
                        pixel_addr <= state_0[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)-160) /320)*80 ]+160;
                    end
                    else if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 3 ) begin
                        pixel_addr <= state_0[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)-240) /320)*80 ]+240;
                    end
                end else if( (h_cnt>>1)+320*(v_cnt>>1) < 51200 ) begin
                    if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 0 ) begin
                        pixel_addr <= state_0[ ( ((h_cnt>>1)+320*(v_cnt>>1))%25600 %320)%80 + ( ((h_cnt>>1)+320*(v_cnt>>1))%25600 /320)*80 ]+25600;
                    end
                    else if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 1 ) begin
                        pixel_addr <= state_0[ ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%25600-80) /320)*80 ]+ 25600 + 80;
                    end
                    else if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 2 ) begin
                        pixel_addr <= state_0[ ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%25600-160) /320)*80 ]+ 25600 + 160;
                    end
                    else if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 3 ) begin
                        pixel_addr <= state_0[ ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%25600-240) /320)*80 ]+ 25600 + 240;
                    end
                end else begin
                    if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 0 ) begin
                        pixel_addr <= state_0[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) /320)*80 ]+51200;
                    end
                    else if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 1 ) begin
                        pixel_addr <= state_0[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200-80) /320)*80 ]+ 51200 + 80;
                    end
                    else if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 2 ) begin
                        pixel_addr <= state_0[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200-160) /320)*80 ]+ 51200 + 160;
                    end
                    else if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 3 ) begin
                        pixel_addr <= state_0[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200-240) /320)*80 ]+ 51200 + 240;
                    end
                end
            end else begin
                
                
                if( (h_cnt>>1)+320*(v_cnt>>1) < 25600 ) begin
                    if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 0 ) begin
                        if(zero == 0) pixel_addr <= state_0[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)) /320)*80 ];
                        else if(zero == 1) pixel_addr <= state_1[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)) /320)*80 ];
                        else if(zero == 2) pixel_addr <= state_2[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)) /320)*80 ];
                        else if(zero == 3) pixel_addr <= state_3[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)) /320)*80 ];
                    end
                    else if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 1 ) begin
                        if(one == 0) pixel_addr <= state_0[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)-80) /320)*80 ]+80;
                        else if(one == 1) pixel_addr <= state_1[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)-80) /320)*80 ]+80;
                        else if(one == 2) pixel_addr <= state_2[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)-80) /320)*80 ]+80;
                        else if(one == 3) pixel_addr <= state_3[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)-80) /320)*80 ]+80;
                    end
                    else if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 2 ) begin
                        if(two == 0) pixel_addr <= state_0[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)-160) /320)*80 ]+160;
                        else if(two == 1) pixel_addr <= state_1[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)-160) /320)*80 ]+160;
                        else if(two == 2) pixel_addr <= state_2[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)-160) /320)*80 ]+160;
                        else if(two == 3) pixel_addr <= state_3[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)-160) /320)*80 ]+160;
                    end
                    else if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 3 ) begin
                        if(three == 0) pixel_addr <= state_0[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)-240) /320)*80 ]+240;
                        else if(three == 1) pixel_addr <= state_1[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)-240) /320)*80 ]+240;
                        else if(three == 2) pixel_addr <= state_2[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)-240) /320)*80 ]+240;
                        else if(three == 3) pixel_addr <= state_3[ (((h_cnt>>1)+320*(v_cnt>>1)) %320)%80 + (((h_cnt>>1)+320*(v_cnt>>1)-240) /320)*80 ]+240;
                    end
                end else if( (h_cnt>>1)+320*(v_cnt>>1) < 51200 ) begin
                    if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 0 ) begin
                        if(four == 0) pixel_addr <= state_0[ ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) /320)*80 ]+25600;
                        else if(four == 1) pixel_addr <= state_1[ ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) /320)*80 ]+25600;
                        else if(four == 2) pixel_addr <= state_2[ ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) /320)*80 ]+25600;
                        else if(four == 3) pixel_addr <= state_3[ ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) /320)*80 ]+25600;
                    end
                    else if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 1 ) begin
                        if(five == 0) pixel_addr <= state_0[ ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%25600-80) /320)*80 ]+ 25600 + 80;
                        else if(five == 1) pixel_addr <= state_1[ ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%25600-80) /320)*80 ]+ 25600 + 80;
                        else if(five == 2) pixel_addr <= state_2[ ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%25600-80) /320)*80 ]+ 25600 + 80;
                        else if(five == 3) pixel_addr <= state_3[ ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%25600-80) /320)*80 ]+ 25600 + 80;
                    end
                    else if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 2 ) begin
                        if(six == 0) pixel_addr <= state_0[ ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%25600-160) /320)*80 ]+ 25600 + 160;
                        else if(six == 1) pixel_addr <= state_1[ ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%25600-160) /320)*80 ]+ 25600 + 160;
                        else if(six == 2) pixel_addr <= state_2[ ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%25600-160) /320)*80 ]+ 25600 + 160;
                        else if(six == 3) pixel_addr <= state_3[ ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%25600-160) /320)*80 ]+ 25600 + 160;
                    end
                    else if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 3 ) begin
                        if(seven == 0) pixel_addr <= state_0[ ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%25600-240) /320)*80 ]+ 25600 + 240;
                        else if(seven == 1) pixel_addr <= state_1[ ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%25600-240) /320)*80 ]+ 25600 + 240;
                        else if(seven == 2) pixel_addr <= state_2[ ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%25600-240) /320)*80 ]+ 25600 + 240;
                        else if(seven == 3) pixel_addr <= state_3[ ( (((h_cnt>>1)+320*(v_cnt>>1))%25600) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%25600-240) /320)*80 ]+ 25600 + 240;
                    end
                end else begin
                    if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 0 ) begin
                        if(eight == 0) pixel_addr <= state_0[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) /320)*80 ]+ 51200;
                        else if(eight == 1) pixel_addr <= state_1[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) /320)*80 ]+ 51200;
                        else if(eight == 2) pixel_addr <= state_2[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) /320)*80 ]+ 51200;
                        else if(eight == 3) pixel_addr <= state_3[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) /320)*80 ]+ 51200;
                    end
                    else if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 1 ) begin
                        if(nine == 0) pixel_addr <= state_0[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200-80) /320)*80 ]+ 51200 + 80;
                        else if(nine == 1) pixel_addr <= state_1[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200-80) /320)*80 ]+ 51200 + 80;
                        else if(nine == 2) pixel_addr <= state_2[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200-80) /320)*80 ]+ 51200 + 80;
                        else if(nine == 3) pixel_addr <= state_3[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200-80) /320)*80 ]+ 51200 + 80;
                    end
                    else if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 2 ) begin
                        if(ten == 0) pixel_addr <= state_0[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200-160) /320)*80 ]+ 51200 + 160;
                        else if(ten == 1) pixel_addr <= state_1[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200-160) /320)*80 ]+ 51200 + 160;
                        else if(ten == 2) pixel_addr <= state_2[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200-160) /320)*80 ]+ 51200 + 160;
                        else if(ten == 3) pixel_addr <= state_3[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200-160) /320)*80 ]+ 51200 + 160;
                    end
                    else if( (((h_cnt>>1)+320*(v_cnt>>1)) %320) / 80 == 3 ) begin
                        if(ele == 0) pixel_addr <= state_0[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200-240) /320)*80 ]+ 51200 + 240;
                        else if(ele == 1) pixel_addr <= state_1[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200-240) /320)*80 ]+ 51200 + 240;
                        else if(ele == 2) pixel_addr <= state_2[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200-240) /320)*80 ]+ 51200 + 240;
                        else if(ele == 3) pixel_addr <= state_3[ ( (((h_cnt>>1)+320*(v_cnt>>1))%51200) %320)%80 + ( (((h_cnt>>1)+320*(v_cnt>>1))%51200-240) /320)*80 ]+ 51200 + 240;
                    end
                end
            end
       
   end
    
    
    
    
    
    
    
    
    
    
    
    
    
    assign {vgaRed, vgaGreen, vgaBlue} = (valid==1'b1) ? pixel : 12'h0;
    assign data = {vgaRed, vgaGreen, vgaBlue};
    blk_mem_gen_0 mem_gen(.addra(pixel_addr), .clka(clk_25MHz), .dina(data), .douta(pixel), .wea(0));
    
endmodule







